CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
176 550 1918 1019
9437202 0
0
6 Title:
5 Name:
0
0
0
5
12 Hex Display~
7 381 85 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3108 0 0
2
43197.7 0
0
12 Hex Display~
7 421 85 0 18 19
10 9 8 7 6 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4299 0 0
2
43197.7 0
0
7 Pulser~
4 169 205 0 10 12
0 11 12 10 13 0 0 10 10 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9672 0 0
2
5.89841e-315 0
0
7 74LS293
154 532 188 0 8 17
0 9 2 6 14 5 4 3 2
0
0 0 4336 0
7 74LS293
-24 -35 25 -27
2 U2
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
5.89841e-315 0
0
7 74LS293
154 346 187 0 8 17
0 9 2 10 9 6 7 8 9
0
0 0 4336 0
7 74LS293
-24 -35 25 -27
2 U1
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
5.89841e-315 0
0
15
1 0 2 0 0 12288 0 1 0 0 9 4
390 109
390 171
437 171
437 245
7 2 3 0 0 12416 0 4 1 0 0 5
564 197
575 197
575 133
384 133
384 109
6 3 4 0 0 12416 0 4 1 0 0 5
564 188
568 188
568 139
378 139
378 109
5 4 5 0 0 8320 0 4 1 0 0 4
564 179
564 145
372 145
372 109
4 0 6 0 0 4224 0 2 0 0 14 4
412 109
412 163
382 163
382 178
6 3 7 0 0 8320 0 5 2 0 0 3
378 187
418 187
418 109
7 2 8 0 0 8320 0 5 2 0 0 3
378 196
424 196
424 109
1 0 9 0 0 4224 0 2 0 0 10 4
430 109
430 210
400 210
400 225
0 2 2 0 0 4224 0 0 5 11 0 4
484 245
291 245
291 187
314 187
0 1 9 0 0 128 0 0 4 15 0 4
378 225
468 225
468 179
500 179
8 2 2 0 0 0 0 4 4 0 0 5
564 206
564 245
483 245
483 188
500 188
0 1 9 0 0 0 0 0 5 15 0 4
308 224
299 224
299 178
314 178
3 3 10 0 0 4224 0 5 3 0 0 2
308 196
193 196
5 3 6 0 0 4224 0 5 4 0 0 4
378 178
442 178
442 197
494 197
4 8 9 0 0 0 0 5 5 0 0 4
308 205
308 225
378 225
378 205
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
