CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 30 100 10
958 88 1917 1018
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
1126 184 1239 281
42991634 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 837 358 0 1 11
0 17
0
0 0 21360 180
2 0V
-7 -16 7 -8
6 Select
-21 -26 21 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6128 0 0
2
43185 0
0
13 Logic Switch~
5 551 143 0 1 11
0 19
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B4
-8 -31 6 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7346 0 0
2
43185 4
0
13 Logic Switch~
5 597 143 0 1 11
0 21
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8577 0 0
2
43185 3
0
13 Logic Switch~
5 691 142 0 1 11
0 23
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3372 0 0
2
43185 2
0
13 Logic Switch~
5 645 142 0 1 11
0 22
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3741 0 0
2
43185 1
0
13 Logic Switch~
5 733 141 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -22 8 -14
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5813 0 0
2
43185 0
0
13 Logic Switch~
5 428 145 0 1 11
0 26
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3213 0 0
2
43185 0
0
13 Logic Switch~
5 340 146 0 1 11
0 28
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3694 0 0
2
43185 1
0
13 Logic Switch~
5 386 146 0 1 11
0 27
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4327 0 0
2
43185 0
0
13 Logic Switch~
5 292 147 0 1 11
0 25
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8800 0 0
2
43185 0
0
13 Logic Switch~
5 246 147 0 1 11
0 20
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3406 0 0
2
43185 0
0
7 Ground~
168 361 486 0 1 3
0 2
0
0 0 53360 180
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6455 0 0
2
43185 0
0
14 Logic Display~
6 689 551 0 1 2
10 12
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9319 0 0
2
43185 0
0
14 Logic Display~
6 689 589 0 1 2
10 13
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S3
-4 -15 10 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3172 0 0
2
43185 0
0
14 Logic Display~
6 689 634 0 1 2
10 14
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
38 0 0
2
43185 0
0
14 Logic Display~
6 689 678 0 1 2
10 15
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
376 0 0
2
43185 0
0
14 Logic Display~
6 690 721 0 1 2
10 16
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S0
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6666 0 0
2
43185 0
0
7 Ground~
168 409 636 0 1 3
0 2
0
0 0 53360 270
0
5 GND10
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9365 0 0
2
43185 0
0
7 Ground~
168 412 670 0 1 3
0 2
0
0 0 53360 270
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3251 0 0
2
43185 0
0
7 Ground~
168 506 679 0 1 3
0 2
0
0 0 53360 90
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5481 0 0
2
43185 0
0
7 74LS151
20 454 698 0 14 29
0 2 33 34 35 36 2 7 6 2
2 2 17 16 37
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
7788 0 0
2
43185 0
0
14 Logic Display~
6 104 415 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Carry
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3273 0 0
2
43185 0
0
7 74LS257
147 454 581 0 14 29
0 17 2 10 2 3 8 4 9 5
2 12 13 14 15
0
0 0 4848 0
7 74LS257
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
3761 0 0
2
43185 0
0
7 Ground~
168 293 432 0 1 3
0 2
0
0 0 53360 90
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3226 0 0
2
43185 0
0
7 Ground~
168 293 396 0 1 3
0 2
0
0 0 53360 90
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4244 0 0
2
43185 0
0
7 74LS283
152 246 424 0 14 29
0 2 2 2 20 2 2 2 19 18
38 39 11 10 40
0
0 0 4848 512
7 74LS283
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
5225 0 0
2
43185 0
0
7 Ground~
168 577 416 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
768 0 0
2
43185 0
0
7 Ground~
168 575 379 0 1 3
0 2
0
0 0 53360 270
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5735 0 0
2
43185 0
0
7 Ground~
168 675 283 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5881 0 0
2
43185 0
0
7 Ground~
168 675 254 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3275 0 0
2
43185 0
0
2 +V
167 693 271 0 1 3
0 32
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4203 0 0
2
43185 0
0
6 74LS85
106 628 398 0 14 29
0 2 2 2 20 2 2 2 19 31
30 29 9 8 7
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
3440 0 0
2
43185 0
0
6 74LS85
106 629 288 0 14 29
0 25 28 27 26 21 22 23 24 2
32 2 31 30 29
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U2
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
9102 0 0
2
43185 0
0
7 Ground~
168 289 341 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5586 0 0
2
43185 0
0
7 74LS283
152 247 297 0 14 29
0 25 28 27 26 21 22 23 24 2
3 4 5 6 18
0
0 0 4848 512
7 74LS283
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
525 0 0
2
43185 0
0
64
0 4 2 0 0 4224 0 0 23 2 0 3
373 494
373 572
422 572
1 2 2 0 0 0 0 12 23 0 0 4
361 494
379 494
379 554
422 554
10 5 3 0 0 8320 0 35 23 0 0 4
215 288
165 288
165 581
422 581
11 7 4 0 0 8320 0 35 23 0 0 4
215 297
173 297
173 599
422 599
12 9 5 0 0 8320 0 35 23 0 0 4
215 306
185 306
185 617
422 617
13 8 6 0 0 8320 0 35 21 0 0 4
215 315
194 315
194 734
422 734
14 7 7 0 0 12416 0 32 21 0 0 6
660 434
671 434
671 493
386 493
386 725
422 725
13 6 8 0 0 12416 0 32 23 0 0 6
660 425
679 425
679 500
393 500
393 590
422 590
12 8 9 0 0 12416 0 32 23 0 0 6
660 416
686 416
686 505
399 505
399 608
422 608
13 3 10 0 0 12416 0 26 23 0 0 4
214 442
202 442
202 563
422 563
12 1 11 0 0 4224 0 26 22 0 0 2
214 433
104 433
11 1 12 0 0 12416 0 23 13 0 0 4
486 563
565 563
565 555
673 555
12 1 13 0 0 12416 0 23 14 0 0 4
486 581
565 581
565 593
673 593
13 1 14 0 0 12416 0 23 15 0 0 4
486 599
549 599
549 638
673 638
14 1 15 0 0 12416 0 23 16 0 0 4
486 617
538 617
538 682
673 682
13 1 16 0 0 4224 0 21 17 0 0 2
486 725
674 725
10 1 2 0 0 0 0 23 18 0 0 2
416 626
416 637
1 0 2 0 0 0 0 19 0 0 19 2
419 671
422 671
6 1 2 0 0 128 0 21 21 0 0 2
422 716
422 671
0 1 2 0 0 0 0 0 20 21 0 4
498 680
504 680
504 680
499 680
10 0 2 0 0 0 0 21 0 0 22 2
486 680
498 680
11 9 2 0 0 0 0 21 21 0 0 4
486 689
498 689
498 671
492 671
12 0 17 0 0 8192 0 21 0 0 24 3
486 698
519 698
519 513
1 1 17 0 0 12416 0 1 23 0 0 6
823 358
692 358
692 513
413 513
413 545
422 545
14 9 18 0 0 16512 0 35 26 0 0 6
215 342
204 342
204 358
313 358
313 469
278 469
8 0 19 0 0 4096 0 26 0 0 35 3
278 451
551 451
551 432
4 0 20 0 0 4096 0 26 0 0 34 3
278 415
462 415
462 398
1 0 2 0 0 0 0 24 0 0 30 2
286 433
286 433
1 0 2 0 0 0 0 25 0 0 32 2
286 397
285 397
6 0 2 0 0 0 0 26 0 0 31 2
278 433
286 433
5 7 2 0 0 0 0 26 26 0 0 4
278 424
286 424
286 442
278 442
2 0 2 0 0 0 0 26 0 0 33 2
278 397
285 397
1 3 2 0 0 0 0 26 26 0 0 4
278 388
285 388
285 406
278 406
1 4 20 0 0 8320 0 11 32 0 0 5
246 159
246 217
462 217
462 398
596 398
1 8 19 0 0 4224 0 2 32 0 0 3
551 155
551 434
596 434
1 0 2 0 0 0 0 27 0 0 37 2
584 417
586 416
6 0 2 0 0 0 0 32 0 0 38 2
596 416
586 416
5 7 2 0 0 128 0 32 32 0 0 4
596 407
586 407
586 425
596 425
1 0 2 0 0 0 0 28 0 0 40 2
582 380
585 380
2 0 2 0 0 0 0 32 0 0 41 2
596 380
585 380
3 1 2 0 0 0 0 32 32 0 0 4
596 389
585 389
585 371
596 371
1 0 21 0 0 12288 0 3 0 0 49 4
597 155
597 193
557 193
557 297
1 0 22 0 0 12288 0 5 0 0 48 4
645 154
645 199
564 199
564 306
1 0 23 0 0 8192 0 4 0 0 47 4
691 154
691 207
572 207
572 315
1 0 24 0 0 8192 0 6 0 0 46 4
733 153
733 215
580 215
580 324
8 8 24 0 0 4224 0 35 33 0 0 2
279 324
597 324
7 7 23 0 0 4224 0 35 33 0 0 2
279 315
597 315
6 6 22 0 0 4224 0 35 33 0 0 2
279 306
597 306
5 5 21 0 0 4224 0 35 33 0 0 2
279 297
597 297
1 0 25 0 0 4096 0 10 0 0 57 2
292 159
292 261
1 0 26 0 0 4096 0 7 0 0 54 2
428 157
428 288
1 0 27 0 0 4096 0 9 0 0 55 2
386 158
386 279
1 0 28 0 0 4096 0 8 0 0 56 2
340 158
340 270
4 4 26 0 0 4224 0 33 35 0 0 2
597 288
279 288
3 3 27 0 0 4224 0 35 33 0 0 2
279 279
597 279
2 2 28 0 0 4224 0 35 33 0 0 2
279 270
597 270
1 1 25 0 0 4224 0 33 35 0 0 2
597 261
279 261
11 14 29 0 0 8320 0 32 33 0 0 4
660 389
680 389
680 324
661 324
13 10 30 0 0 8320 0 33 32 0 0 4
661 315
674 315
674 380
660 380
9 12 31 0 0 8320 0 32 33 0 0 4
660 371
666 371
666 306
661 306
11 1 2 0 0 0 0 33 29 0 0 3
661 279
661 284
668 284
1 9 2 0 0 0 0 30 33 0 0 3
668 255
661 255
661 261
1 10 32 0 0 4224 0 31 33 0 0 2
681 270
661 270
1 9 2 0 0 0 0 34 35 0 0 4
282 342
291 342
291 342
279 342
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
