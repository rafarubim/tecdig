CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 20 30 100 10
1137 88 1917 1018
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
1305 184 1418 281
42991634 0
0
6 Title:
5 Name:
0
0
0
41
13 Logic Switch~
5 591 156 0 1 11
0 36
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5435 0 0
2
43192 0
0
13 Logic Switch~
5 629 156 0 1 11
0 41
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3446 0 0
2
43192 0
0
13 Logic Switch~
5 664 157 0 1 11
0 40
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3914 0 0
2
43192 0
0
13 Logic Switch~
5 699 158 0 1 11
0 39
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3948 0 0
2
43192 0
0
13 Logic Switch~
5 733 158 0 1 11
0 38
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3901 0 0
2
43192 0
0
13 Logic Switch~
5 369 157 0 1 11
0 37
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A4
-6 -32 8 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6295 0 0
2
43192 0
0
13 Logic Switch~
5 405 158 0 1 11
0 45
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A3
-6 -32 8 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
332 0 0
2
43192 0
0
13 Logic Switch~
5 439 160 0 1 11
0 44
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A2
-6 -32 8 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9737 0 0
2
43192 0
0
13 Logic Switch~
5 474 160 0 1 11
0 43
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A1
-6 -32 8 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9910 0 0
2
43192 0
0
13 Logic Switch~
5 511 160 0 1 11
0 42
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A0
-6 -32 8 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3834 0 0
2
43192 0
0
7 Ground~
168 662 794 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3138 0 0
2
43192 0
0
14 Logic Display~
6 844 768 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 CONV
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5409 0 0
2
43192 0
0
2 +V
167 665 696 0 1 3
0 6
0
0 0 53744 90
2 5V
-7 -15 7 -7
0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
983 0 0
2
43192 0
0
7 Ground~
168 669 666 0 1 3
0 2
0
0 0 53360 270
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6652 0 0
2
43192 0
0
7 Ground~
168 782 639 0 1 3
0 2
0
0 0 53360 90
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4281 0 0
2
43192 0
0
6 74LS85
106 731 768 0 14 29
0 2 2 5 4 2 2 2 6 7
8 9 3 47 48
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U7
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
6847 0 0
2
43192 0
0
6 74LS85
106 731 658 0 14 29
0 13 12 11 10 2 2 6 6 2
2 2 7 8 9
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U6
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
6543 0 0
2
43192 0
0
7 Ground~
168 386 720 0 1 3
0 2
0
0 0 53360 270
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7168 0 0
2
43192 0
0
12 Hex Display~
7 607 684 0 16 19
10 19 20 21 22 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3828 0 0
2
43192 0
0
12 Hex Display~
7 565 684 0 16 19
10 15 16 17 18 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
955 0 0
2
43192 0
0
7 Ground~
168 381 832 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7782 0 0
2
43192 0
0
9 Inverter~
13 411 545 0 2 22
0 24 14
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U5A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
824 0 0
2
43192 0
0
7 74LS283
152 432 806 0 14 29
0 2 2 5 4 2 2 2 2 23
18 17 16 15 49
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 S4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
6983 0 0
2
43192 0
0
7 74LS283
152 434 676 0 14 29
0 13 12 11 10 2 14 14 2 2
22 21 20 19 23
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 S3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
3185 0 0
2
43192 0
0
8 2-In OR~
219 459 545 0 3 22
0 25 5 24
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U4A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4213 0 0
2
43192 0
0
9 Inverter~
13 760 554 0 2 22
0 26 25
0
0 0 624 180
6 74LS04
-21 -19 21 -11
2 NF
-1 -20 13 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
9765 0 0
2
43192 0
0
8 4-In OR~
219 808 519 0 5 22
0 27 28 29 30 26
0
0 0 624 270
4 4072
-14 -24 14 -16
3 U3A
26 -5 47 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
8986 0 0
2
43192 0
0
9 4-In AND~
219 765 428 0 5 22
0 4 33 32 34 29
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
3273 0 0
2
43192 0
0
9 4-In AND~
219 766 481 0 5 22
0 4 33 32 31 30
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 3 0
1 U
5636 0 0
2
43192 0
0
9 3-In AND~
219 765 378 0 4 22
0 35 13 12 28
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 2 0
1 U
327 0 0
2
43192 0
0
9 3-In AND~
219 764 331 0 4 22
0 35 13 11 27
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
9233 0 0
2
43192 0
0
9 Inverter~
13 719 297 0 2 22
0 10 31
0
0 0 624 270
6 74LS04
-21 -19 21 -11
2 NE
19 -8 33 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3875 0 0
2
43192 0
0
9 Inverter~
13 668 299 0 2 22
0 11 34
0
0 0 624 270
6 74LS04
-21 -19 21 -11
2 ND
19 -8 33 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9991 0 0
2
43192 0
0
9 Inverter~
13 617 300 0 2 22
0 12 32
0
0 0 624 270
6 74LS04
-21 -19 21 -11
2 NC
19 -8 33 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3221 0 0
2
43192 0
0
9 Inverter~
13 565 301 0 2 22
0 13 33
0
0 0 624 270
6 74LS04
-21 -19 21 -11
2 NB
19 -8 33 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8874 0 0
2
43192 0
0
9 Inverter~
13 512 301 0 2 22
0 4 35
0
0 0 624 270
6 74LS04
-21 -19 21 -11
2 NA
19 -8 33 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7400 0 0
2
43192 0
0
7 Ground~
168 372 455 0 1 3
0 2
0
0 0 53360 270
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3623 0 0
2
43192 0
0
7 Ground~
168 372 419 0 1 3
0 2
0
0 0 53360 270
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3311 0 0
2
43192 0
0
7 Ground~
168 392 357 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5736 0 0
2
43192 0
0
7 74LS283
152 431 447 0 14 29
0 2 2 2 37 2 2 2 36 46
50 51 5 4 52
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 S2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
3143 0 0
2
43192 0
0
7 74LS283
152 430 313 0 14 29
0 45 44 43 42 41 40 39 38 2
13 12 11 10 46
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 S1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
5835 0 0
2
43192 0
0
99
0 1 2 0 0 4096 0 0 11 14 0 2
690 795
669 795
11 0 2 0 0 0 0 17 0 0 3 3
763 649
770 649
770 640
9 0 2 0 0 0 0 17 0 0 19 3
763 631
770 631
770 640
12 1 3 0 0 4224 0 16 12 0 0 2
763 786
844 786
0 4 4 0 0 8192 0 0 16 38 0 5
501 565
501 634
642 634
642 768
699 768
0 3 5 0 0 8192 0 0 16 37 0 5
491 575
491 627
648 627
648 759
699 759
0 1 2 0 0 0 0 0 16 8 0 3
690 750
690 741
699 741
2 0 2 0 0 8320 0 16 0 0 15 3
699 750
690 750
690 777
8 1 6 0 0 8320 0 16 13 0 0 3
699 804
676 804
676 694
1 0 6 0 0 0 0 13 0 0 11 2
676 694
676 694
7 8 6 0 0 0 0 17 17 0 0 4
699 685
676 685
676 694
699 694
6 1 2 0 0 0 0 17 14 0 0 3
699 676
676 676
676 667
1 5 2 0 0 0 0 14 17 0 0 2
676 667
699 667
7 0 2 0 0 0 0 16 0 0 15 3
699 795
690 795
690 786
6 5 2 0 0 0 0 16 16 0 0 4
699 786
690 786
690 777
699 777
12 9 7 0 0 8320 0 17 16 0 0 4
763 676
778 676
778 741
763 741
13 10 8 0 0 8320 0 17 16 0 0 4
763 685
773 685
773 750
763 750
14 11 9 0 0 8320 0 17 16 0 0 4
763 694
768 694
768 759
763 759
10 1 2 0 0 0 0 17 15 0 0 2
763 640
775 640
0 4 10 0 0 4096 0 0 17 82 0 3
681 582
681 658
699 658
0 3 11 0 0 8192 0 0 17 83 0 5
656 592
656 622
687 622
687 649
699 649
0 2 12 0 0 8192 0 0 17 84 0 5
603 598
603 616
693 616
693 640
699 640
0 1 13 0 0 4096 0 0 17 85 0 3
551 610
699 610
699 631
8 0 2 0 0 0 0 24 0 0 25 2
402 703
393 703
5 1 2 0 0 8192 0 24 18 0 0 3
402 676
393 676
393 721
9 1 2 0 0 0 0 24 18 0 0 2
402 721
393 721
7 0 14 0 0 4096 0 24 0 0 55 3
402 694
372 694
372 685
0 1 10 0 0 0 0 0 32 82 0 3
705 270
722 270
722 279
0 1 11 0 0 0 0 0 33 83 0 3
656 262
671 262
671 281
0 1 12 0 0 0 0 0 34 84 0 3
603 255
620 255
620 282
0 1 13 0 0 0 0 0 35 85 0 3
549 249
568 249
568 283
2 0 2 0 0 0 0 23 0 0 52 2
400 779
388 779
5 0 2 0 0 0 0 23 0 0 52 2
400 806
388 806
6 0 2 0 0 0 0 23 0 0 52 2
400 815
388 815
7 0 2 0 0 0 0 23 0 0 52 2
400 824
388 824
2 0 5 0 0 0 0 25 0 0 37 2
478 536
491 536
12 3 5 0 0 16512 0 40 23 0 0 6
463 456
491 456
491 575
365 575
365 788
400 788
0 4 4 0 0 12288 0 0 23 67 0 5
501 468
501 567
357 567
357 797
400 797
0 13 4 0 0 0 0 0 40 71 0 4
501 243
484 243
484 465
463 465
0 7 2 0 0 0 0 0 40 41 0 3
393 456
393 465
399 465
5 0 2 0 0 0 0 40 0 0 88 3
399 447
393 447
393 456
1 0 2 0 0 0 0 40 0 0 43 3
399 411
393 411
393 420
3 0 2 0 0 0 0 40 0 0 89 3
399 429
393 429
393 420
13 1 15 0 0 8320 0 23 20 0 0 3
464 824
574 824
574 708
12 2 16 0 0 8320 0 23 20 0 0 3
464 815
568 815
568 708
11 3 17 0 0 4224 0 23 20 0 0 3
464 806
562 806
562 708
10 4 18 0 0 4224 0 23 20 0 0 3
464 797
556 797
556 708
13 1 19 0 0 12416 0 24 19 0 0 5
466 694
525 694
525 726
616 726
616 708
12 2 20 0 0 12416 0 24 19 0 0 5
466 685
531 685
531 721
610 721
610 708
11 3 21 0 0 4224 0 24 19 0 0 5
466 676
536 676
536 716
604 716
604 708
10 4 22 0 0 4224 0 24 19 0 0 5
466 667
541 667
541 711
598 711
598 708
1 1 2 0 0 4224 0 21 23 0 0 3
388 833
388 770
400 770
8 1 2 0 0 0 0 23 21 0 0 2
400 833
388 833
14 9 23 0 0 16512 0 24 23 0 0 6
466 721
469 721
469 739
394 739
394 851
400 851
2 6 14 0 0 8320 0 22 24 0 0 4
396 545
372 545
372 685
402 685
1 3 24 0 0 0 0 22 25 0 0 2
432 545
432 545
1 2 25 0 0 4224 0 25 26 0 0 2
478 554
745 554
1 5 26 0 0 4224 0 26 27 0 0 3
781 554
811 554
811 549
4 1 27 0 0 8320 0 31 27 0 0 3
785 331
824 331
824 499
4 2 28 0 0 8320 0 30 27 0 0 3
786 378
815 378
815 499
5 3 29 0 0 8320 0 28 27 0 0 3
786 428
806 428
806 499
5 4 30 0 0 8320 0 29 27 0 0 3
787 481
797 481
797 499
4 0 31 0 0 4096 0 29 0 0 64 2
742 495
722 495
2 0 31 0 0 4224 0 32 0 0 0 2
722 315
722 507
3 0 32 0 0 4096 0 29 0 0 79 2
742 486
620 486
2 0 33 0 0 4096 0 29 0 0 80 2
742 477
568 477
1 0 4 0 0 4224 0 29 0 0 71 3
742 468
501 468
501 415
4 0 34 0 0 4096 0 28 0 0 78 2
741 442
671 442
3 0 32 0 0 0 0 28 0 0 79 2
741 433
620 433
2 0 33 0 0 0 0 28 0 0 80 2
741 424
568 424
1 1 4 0 0 0 0 28 36 0 0 5
741 415
501 415
501 243
515 243
515 283
3 0 12 0 0 4096 0 30 0 0 84 2
741 387
603 387
2 0 13 0 0 4096 0 30 0 0 85 2
741 378
551 378
1 0 35 0 0 4224 0 30 0 0 81 2
741 369
515 369
3 0 11 0 0 4096 0 31 0 0 83 2
740 340
656 340
2 0 13 0 0 0 0 31 0 0 85 2
740 331
551 331
1 0 35 0 0 0 0 31 0 0 81 2
740 322
515 322
2 0 34 0 0 4224 0 33 0 0 0 2
671 317
671 507
2 0 32 0 0 4224 0 34 0 0 0 2
620 318
620 507
2 0 33 0 0 4224 0 35 0 0 0 2
568 319
568 507
2 0 35 0 0 0 0 36 0 0 0 2
515 319
515 507
13 4 10 0 0 20608 0 41 24 0 0 8
462 331
479 331
479 270
705 270
705 582
380 582
380 667
402 667
12 3 11 0 0 16512 0 41 24 0 0 8
462 322
475 322
475 262
656 262
656 592
388 592
388 658
402 658
11 2 12 0 0 16512 0 41 24 0 0 8
462 313
468 313
468 255
603 255
603 600
395 600
395 649
402 649
10 1 13 0 0 12416 0 41 24 0 0 6
462 304
462 249
551 249
551 610
402 610
402 640
1 8 36 0 0 12416 0 1 40 0 0 5
591 168
591 195
340 195
340 474
399 474
1 4 37 0 0 12416 0 6 40 0 0 5
369 169
369 202
348 202
348 438
399 438
1 6 2 0 0 0 0 37 40 0 0 2
379 456
399 456
1 2 2 0 0 0 0 38 40 0 0 2
379 420
399 420
1 8 38 0 0 8320 0 5 41 0 0 5
733 170
733 208
356 208
356 340
398 340
1 7 39 0 0 8320 0 4 41 0 0 5
699 170
699 216
363 216
363 331
398 331
1 6 40 0 0 8320 0 3 41 0 0 5
664 169
664 223
370 223
370 322
398 322
1 5 41 0 0 8320 0 2 41 0 0 5
629 168
629 229
376 229
376 313
398 313
1 4 42 0 0 8320 0 10 41 0 0 5
511 172
511 235
382 235
382 304
398 304
1 3 43 0 0 8320 0 9 41 0 0 5
474 172
474 241
387 241
387 295
398 295
1 2 44 0 0 4224 0 8 41 0 0 5
439 172
439 247
393 247
393 286
398 286
1 1 45 0 0 4224 0 7 41 0 0 4
405 170
405 251
398 251
398 277
14 9 46 0 0 16512 0 41 40 0 0 6
462 358
477 358
477 377
389 377
389 492
399 492
1 9 2 0 0 0 0 39 41 0 0 2
399 358
398 358
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
