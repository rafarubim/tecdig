CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
1180 88 1917 1018
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
1348 184 1461 281
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 268 629 0 1 11
0 16
0
0 0 21360 90
2 0V
11 0 25 8
1 E
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4139 0 0
2
43178.2 0
0
13 Logic Switch~
5 214 628 0 1 11
0 17
0
0 0 21360 90
2 0V
11 0 25 8
1 D
13 -10 20 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6435 0 0
2
43178.2 0
0
13 Logic Switch~
5 159 627 0 1 11
0 18
0
0 0 21360 90
2 0V
11 0 25 8
1 C
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5283 0 0
2
43178.2 0
0
13 Logic Switch~
5 106 626 0 1 11
0 19
0
0 0 21360 90
2 0V
11 0 25 8
1 B
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6874 0 0
2
43178.2 0
0
13 Logic Switch~
5 60 624 0 1 11
0 20
0
0 0 21360 90
2 0V
11 0 25 8
1 A
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5305 0 0
2
43178.2 0
0
5 4049~
219 255 453 0 2 22
0 16 21
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4E
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
34 0 0
2
43178.2 0
0
5 4049~
219 200 481 0 2 22
0 17 22
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4D
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
969 0 0
2
43178.2 0
0
5 4049~
219 147 443 0 2 22
0 18 23
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4C
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
8402 0 0
2
43178.2 0
0
5 4049~
219 95 482 0 2 22
0 19 24
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4B
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
3751 0 0
2
43178.2 0
0
5 4049~
219 60 438 0 2 22
0 20 25
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4A
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
4292 0 0
2
43178.2 0
0
7 Ground~
168 720 418 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6118 0 0
2
43178.2 0
0
4 LED~
171 666 418 0 2 2
10 3 2
0
0 0 864 90
4 LED1
-12 -21 16 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
34 0 0
2
43178.2 0
0
8 2-In OR~
219 608 420 0 3 22
0 4 5 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6357 0 0
2
43178.2 0
0
8 2-In OR~
219 544 525 0 3 22
0 6 7 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
319 0 0
2
43178.2 0
0
8 2-In OR~
219 541 312 0 3 22
0 9 8 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3976 0 0
2
43178.2 0
0
8 2-In OR~
219 477 472 0 3 22
0 11 10 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7634 0 0
2
43178.2 0
0
8 2-In OR~
219 482 367 0 3 22
0 13 12 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
523 0 0
2
43178.2 0
0
8 2-In OR~
219 485 256 0 3 22
0 15 14 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6748 0 0
2
43178.2 0
0
9 3-In AND~
219 402 543 0 4 22
0 20 19 17 7
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 3 0
1 U
6901 0 0
2
43178.1 0
0
9 3-In AND~
219 402 496 0 4 22
0 20 19 18 10
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 3 0
1 U
842 0 0
2
43178.1 0
0
9 4-In AND~
219 403 449 0 5 22
0 20 24 23 16 11
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
3277 0 0
2
43178.1 0
0
9 3-In AND~
219 402 396 0 4 22
0 19 23 17 12
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
4212 0 0
2
43178.1 0
0
9 4-In AND~
219 402 341 0 5 22
0 25 23 17 21 13
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
4720 0 0
2
43178.1 0
0
9 4-In AND~
219 401 288 0 5 22
0 25 19 22 16 14
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U1B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
5551 0 0
2
43178.1 0
0
9 4-In AND~
219 401 236 0 5 22
0 25 24 23 22 15
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U1A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 1 0
1 U
6986 0 0
2
43178.1 0
0
46
2 1 2 0 0 4224 0 12 11 0 0 2
679 419
713 419
3 1 3 0 0 8320 0 13 12 0 0 3
641 420
641 419
659 419
1 3 4 0 0 8320 0 13 15 0 0 4
595 411
582 411
582 312
574 312
3 2 5 0 0 8320 0 14 13 0 0 4
577 525
587 525
587 429
595 429
1 3 6 0 0 8320 0 14 16 0 0 4
531 516
518 516
518 472
510 472
4 2 7 0 0 4224 0 19 14 0 0 4
423 543
523 543
523 534
531 534
3 2 8 0 0 8320 0 17 15 0 0 4
515 367
520 367
520 321
528 321
3 1 9 0 0 8320 0 18 15 0 0 4
518 256
522 256
522 303
528 303
4 2 10 0 0 4224 0 20 16 0 0 4
423 496
456 496
456 481
464 481
5 1 11 0 0 4224 0 21 16 0 0 4
424 449
456 449
456 463
464 463
4 2 12 0 0 4224 0 22 17 0 0 4
423 396
461 396
461 376
469 376
5 1 13 0 0 4224 0 23 17 0 0 4
423 341
461 341
461 358
469 358
5 2 14 0 0 4224 0 24 18 0 0 4
422 288
464 288
464 265
472 265
5 1 15 0 0 4224 0 25 18 0 0 4
422 236
464 236
464 247
472 247
4 0 16 0 0 4096 0 21 0 0 16 2
379 463
325 463
0 4 16 0 0 16512 0 0 24 42 0 6
258 571
269 571
269 572
325 572
325 302
377 302
3 0 17 0 0 4096 0 19 0 0 19 3
378 552
280 552
280 535
3 0 17 0 0 0 0 22 0 0 19 2
378 405
280 405
0 3 17 0 0 12416 0 0 23 43 0 5
203 536
203 535
280 535
280 346
378 346
0 0 18 0 0 8192 0 0 0 21 44 3
165 524
165 525
151 525
0 3 18 0 0 4224 0 0 20 0 0 4
159 524
313 524
313 505
378 505
2 0 19 0 0 4096 0 19 0 0 26 5
378 543
315 543
315 542
305 542
305 514
0 2 19 0 0 4096 0 0 20 26 0 4
305 497
370 497
370 496
378 496
0 1 19 0 0 4096 0 0 22 26 0 2
305 387
378 387
0 0 19 0 0 0 0 0 0 26 45 3
106 514
106 515
98 515
0 2 19 0 0 8320 0 0 24 0 0 4
103 514
305 514
305 284
377 284
1 0 20 0 0 4096 0 19 0 0 29 3
378 534
298 534
298 506
1 0 20 0 0 0 0 20 0 0 29 2
378 487
298 487
0 1 20 0 0 4224 0 0 21 46 0 4
63 506
298 506
298 436
379 436
2 4 21 0 0 16512 0 6 23 0 0 5
258 435
258 427
259 427
259 355
378 355
3 0 22 0 0 4096 0 24 0 0 32 4
377 293
208 293
208 294
203 294
2 4 22 0 0 4224 0 7 25 0 0 3
203 463
203 250
377 250
3 0 23 0 0 16384 0 21 0 0 34 5
379 454
372 454
372 453
333 453
333 396
2 0 23 0 0 4224 0 22 0 0 36 2
378 396
151 396
2 0 23 0 0 0 0 23 0 0 36 2
378 337
151 337
2 3 23 0 0 0 0 8 25 0 0 4
150 425
151 425
151 241
377 241
2 0 24 0 0 20480 0 21 0 0 38 6
379 445
368 445
368 446
292 446
292 412
98 412
2 2 24 0 0 8320 0 9 25 0 0 3
98 464
98 232
377 232
1 0 25 0 0 4224 0 23 0 0 41 2
378 328
62 328
1 0 25 0 0 0 0 24 0 0 41 2
377 275
62 275
2 1 25 0 0 0 0 10 25 0 0 5
63 420
63 390
62 390
62 223
377 223
1 1 16 0 0 0 0 6 1 0 0 4
258 471
258 609
269 609
269 616
1 1 17 0 0 0 0 7 2 0 0 4
203 499
203 608
215 608
215 615
1 1 18 0 0 0 0 8 3 0 0 5
150 461
151 461
151 607
160 607
160 614
1 1 19 0 0 0 0 9 4 0 0 4
98 500
98 606
107 606
107 613
1 1 20 0 0 0 0 10 5 0 0 4
63 456
63 604
61 604
61 611
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
