CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
897 88 1437 838
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
1065 184 1178 281
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 276 66 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43192 0
0
13 Logic Switch~
5 84 600 0 1 11
0 5
0
0 0 21360 90
2 0V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43192 0
0
13 Logic Switch~
5 50 600 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43192 0
0
13 Logic Switch~
5 86 476 0 1 11
0 7
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43192 0
0
13 Logic Switch~
5 49 475 0 1 11
0 4
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43192 0
0
13 Logic Switch~
5 86 342 0 1 11
0 8
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43192 0
0
13 Logic Switch~
5 50 342 0 1 11
0 9
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43192 0
0
13 Logic Switch~
5 85 214 0 1 11
0 10
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43192 0
0
13 Logic Switch~
5 49 214 0 1 11
0 11
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4747 0 0
2
43192 0
0
13 Logic Switch~
5 404 693 0 1 11
0 13
0
0 0 21360 90
2 0V
11 0 25 8
2 S2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43192 0
0
13 Logic Switch~
5 346 692 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
2 S1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
43192 0
0
13 Logic Switch~
5 288 691 0 1 11
0 15
0
0 0 21360 90
2 0V
11 0 25 8
2 S0
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
43192 0
0
14 Logic Display~
6 499 357 0 1 2
10 12
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43192 0
0
7 Ground~
168 208 633 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4597 0 0
2
43192 0
0
7 Ground~
168 41 631 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3835 0 0
2
43192 0
0
7 74LS151
20 399 335 0 14 29
0 2 2 2 2 2 2 16 17 3
2 2 13 12 22
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
3670 0 0
2
43192 0
0
7 74LS151
20 278 469 0 14 29
0 2 2 2 2 2 2 19 18 3
2 2 14 17 23
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
5616 0 0
2
43192 0
0
7 74LS151
20 277 218 0 14 29
0 2 2 2 2 2 2 21 20 3
2 2 14 16 24
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
9323 0 0
2
43192 0
0
7 74LS151
20 135 537 0 14 29
0 2 2 2 2 2 2 6 5 3
2 2 15 18 25
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
317 0 0
2
43192 0
0
7 74LS151
20 134 405 0 14 29
0 2 2 2 2 2 2 4 7 3
2 2 15 19 26
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
3108 0 0
2
43192 0
0
7 74LS151
20 132 277 0 14 29
0 2 2 2 2 2 2 9 8 3
2 2 15 20 27
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
4299 0 0
2
43192 0
0
7 74LS151
20 131 150 0 14 29
0 2 2 2 2 2 2 11 10 3
2 2 15 21 28
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
9672 0 0
2
43192 0
0
85
9 0 3 0 0 8192 0 21 0 0 3 3
170 250
173 250
173 242
0 9 3 0 0 0 0 0 20 3 0 3
173 381
172 381
172 378
9 0 3 0 0 4224 0 19 0 0 7 2
173 510
173 123
9 9 3 0 0 0 0 17 18 0 0 3
316 442
315 442
315 191
9 0 3 0 0 0 0 16 0 0 6 3
437 308
437 123
315 123
9 0 3 0 0 0 0 18 0 0 7 3
315 191
315 123
275 123
9 1 3 0 0 0 0 22 1 0 0 3
169 123
276 123
276 78
1 7 4 0 0 8320 0 5 20 0 0 3
50 462
50 432
102 432
1 8 5 0 0 8320 0 2 19 0 0 3
85 587
85 573
103 573
1 7 6 0 0 8320 0 3 19 0 0 3
51 587
51 564
103 564
1 8 7 0 0 4224 0 4 20 0 0 3
87 463
87 441
102 441
1 8 8 0 0 4224 0 6 21 0 0 3
87 329
87 313
100 313
1 7 9 0 0 8320 0 7 21 0 0 3
51 329
51 304
100 304
1 8 10 0 0 4224 0 8 22 0 0 3
86 201
86 186
99 186
1 7 11 0 0 8320 0 9 22 0 0 3
50 201
50 177
99 177
13 1 12 0 0 8320 0 16 13 0 0 3
431 362
431 361
483 361
1 12 13 0 0 12416 0 10 16 0 0 5
405 680
405 601
466 601
466 335
431 335
12 0 14 0 0 4096 0 17 0 0 19 2
310 469
347 469
1 12 14 0 0 4224 0 11 18 0 0 3
347 679
347 218
309 218
12 0 15 0 0 4096 0 19 0 0 23 2
167 537
186 537
12 0 15 0 0 4096 0 20 0 0 23 2
166 405
186 405
12 0 15 0 0 4096 0 21 0 0 23 2
164 277
186 277
1 12 15 0 0 12416 0 12 22 0 0 5
289 678
289 601
186 601
186 150
163 150
10 0 2 0 0 4096 0 16 0 0 25 2
431 317
466 317
11 0 2 0 0 12288 0 16 0 0 28 4
431 326
466 326
466 209
328 209
10 0 2 0 0 0 0 17 0 0 27 2
310 451
328 451
11 0 2 0 0 0 0 17 0 0 30 3
310 460
328 460
328 353
11 0 2 0 0 0 0 18 0 0 29 2
309 209
328 209
10 0 2 0 0 0 0 18 0 0 35 3
309 200
328 200
328 308
6 0 2 0 0 4096 0 16 0 0 61 2
367 353
208 353
5 0 2 0 0 0 0 16 0 0 61 2
367 344
208 344
4 0 2 0 0 0 0 16 0 0 61 2
367 335
208 335
3 0 2 0 0 0 0 16 0 0 61 2
367 326
208 326
2 0 2 0 0 0 0 16 0 0 61 2
367 317
208 317
1 0 2 0 0 0 0 16 0 0 61 2
367 308
208 308
13 7 16 0 0 8320 0 18 16 0 0 4
309 245
340 245
340 362
367 362
13 8 17 0 0 8320 0 17 16 0 0 4
310 496
340 496
340 371
367 371
6 0 2 0 0 0 0 17 0 0 61 2
246 487
208 487
5 0 2 0 0 0 0 17 0 0 61 2
246 478
208 478
4 0 2 0 0 0 0 17 0 0 61 2
246 469
208 469
3 0 2 0 0 0 0 17 0 0 61 2
246 460
208 460
2 0 2 0 0 0 0 17 0 0 61 2
246 451
208 451
1 0 2 0 0 0 0 17 0 0 61 2
246 442
208 442
6 0 2 0 0 0 0 18 0 0 61 2
245 236
208 236
5 0 2 0 0 0 0 18 0 0 61 2
245 227
208 227
4 0 2 0 0 0 0 18 0 0 61 2
245 218
208 218
3 0 2 0 0 0 0 18 0 0 61 2
245 209
208 209
2 0 2 0 0 0 0 18 0 0 61 2
245 200
208 200
1 0 2 0 0 0 0 18 0 0 61 2
245 191
208 191
13 8 18 0 0 8320 0 19 17 0 0 4
167 564
223 564
223 505
246 505
13 7 19 0 0 8320 0 20 17 0 0 4
166 432
223 432
223 496
246 496
13 8 20 0 0 4224 0 21 18 0 0 4
164 304
223 304
223 254
245 254
13 7 21 0 0 8320 0 22 18 0 0 4
163 177
223 177
223 245
245 245
11 0 2 0 0 0 0 19 0 0 61 2
167 528
208 528
10 0 2 0 0 0 0 19 0 0 61 2
167 519
208 519
11 0 2 0 0 0 0 20 0 0 61 2
166 396
208 396
10 0 2 0 0 0 0 20 0 0 61 2
166 387
208 387
11 0 2 0 0 0 0 21 0 0 61 2
164 268
208 268
10 0 2 0 0 0 0 21 0 0 61 2
164 259
208 259
11 0 2 0 0 0 0 22 0 0 61 2
163 141
208 141
1 10 2 0 0 4096 0 14 22 0 0 3
208 627
208 132
163 132
6 0 2 0 0 0 0 19 0 0 85 2
103 555
41 555
5 0 2 0 0 0 0 19 0 0 85 2
103 546
41 546
4 0 2 0 0 0 0 19 0 0 85 2
103 537
41 537
3 0 2 0 0 0 0 19 0 0 85 2
103 528
41 528
2 0 2 0 0 0 0 19 0 0 85 2
103 519
41 519
1 0 2 0 0 0 0 19 0 0 85 2
103 510
41 510
6 0 2 0 0 0 0 20 0 0 85 2
102 423
41 423
5 0 2 0 0 0 0 20 0 0 85 2
102 414
41 414
4 0 2 0 0 0 0 20 0 0 85 2
102 405
41 405
3 0 2 0 0 0 0 20 0 0 85 2
102 396
41 396
2 0 2 0 0 0 0 20 0 0 85 2
102 387
41 387
1 0 2 0 0 0 0 20 0 0 85 2
102 378
41 378
6 0 2 0 0 0 0 21 0 0 85 2
100 295
41 295
5 0 2 0 0 0 0 21 0 0 85 2
100 286
41 286
4 0 2 0 0 0 0 21 0 0 85 2
100 277
41 277
3 0 2 0 0 0 0 21 0 0 85 2
100 268
41 268
2 0 2 0 0 0 0 21 0 0 85 2
100 259
41 259
1 0 2 0 0 0 0 21 0 0 85 2
100 250
41 250
6 0 2 0 0 0 0 22 0 0 85 2
99 168
41 168
5 0 2 0 0 0 0 22 0 0 85 2
99 159
41 159
4 0 2 0 0 0 0 22 0 0 85 2
99 150
41 150
3 0 2 0 0 0 0 22 0 0 85 2
99 141
41 141
2 0 2 0 0 0 0 22 0 0 85 2
99 132
41 132
1 1 2 0 0 4224 0 15 22 0 0 3
41 625
41 123
99 123
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
