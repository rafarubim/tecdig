CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 100 10
647 129 1551 1059
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
815 225 928 322
9437202 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 204 171 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
4 MODO
-13 -31 15 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
828 0 0
2
43232.7 0
0
9 2-In AND~
219 484 595 0 3 22
0 4 5 6
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U7C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6187 0 0
2
43232.8 0
0
9 2-In NOR~
219 451 538 0 3 22
0 7 8 5
0
0 0 112 270
6 74LS02
-21 -24 21 -16
3 U4A
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7107 0 0
2
43232.8 0
0
2 +V
167 528 523 0 1 3
0 9
0
0 0 53360 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6433 0 0
2
43232.8 0
0
5 7425~
219 502 539 0 6 22
0 21 22 23 24 9 4
0
0 0 112 270
4 7425
-14 -24 14 -16
4 U10A
-6 19 22 27
0
15 DVCC=14;DGND=7;
69 %D [%14bi %7bi %1i %2i %3i %4i %5i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 5 4 2 1 3 6 5 4 2
1 3 6 9 10 12 13 11 8 0
0 6 0
65 0 0 0 2 1 6 0
1 U
8559 0 0
2
43232.8 0
0
9 2-In AND~
219 551 547 0 3 22
0 22 3 26
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U7B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3674 0 0
2
43232.8 0
0
2 +V
167 639 205 0 1 3
0 10
0
0 0 53360 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5697 0 0
2
43232.8 0
0
7 Ground~
168 617 205 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3805 0 0
2
43232.8 0
0
7 Ground~
168 652 355 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5219 0 0
2
43232.8 0
0
7 Ground~
168 312 543 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3795 0 0
2
43232.8 0
0
7 74LS157
122 695 295 0 14 29
0 11 2 2 2 2 10 2 2 2
2 13 14 15 16
0
0 0 4336 0
7 74LS157
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
3637 0 0
2
43232.8 0
0
2 +V
167 268 434 0 1 3
0 12
0
0 0 53360 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3226 0 0
2
43232.8 0
0
7 Ground~
168 250 433 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6966 0 0
2
43232.8 0
0
7 74LS157
122 352 476 0 14 29
0 11 2 2 2 12 12 12 12 12
2 20 19 18 17
0
0 0 4336 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
9796 0 0
2
43232.8 0
0
8 2-In OR~
219 422 632 0 3 22
0 26 6 25
0
0 0 112 180
6 74LS32
-21 -24 21 -16
3 U5A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5952 0 0
2
43232.7 0
0
9 Inverter~
13 333 574 0 2 22
0 25 27
0
0 0 112 180
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3649 0 0
2
43232.7 0
0
12 Hex Display~
7 500 423 0 16 19
10 21 22 23 24 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3716 0 0
2
43232.7 0
0
12 Hex Display~
7 540 423 0 18 19
10 7 28 3 8 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4797 0 0
2
43232.7 0
0
7 74LS190
134 557 321 0 14 29
0 30 29 27 11 13 14 15 16 32
33 24 23 22 21
0
0 0 4336 0
7 74LS190
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
4681 0 0
2
43232.7 0
0
9 Inverter~
13 456 315 0 2 22
0 31 30
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9730 0 0
2
43232.7 0
0
7 Ground~
168 324 266 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9874 0 0
2
43232.7 0
0
7 Pulser~
4 154 306 0 10 12
0 34 35 29 36 0 0 10 10 7
7
0
0 0 4144 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
364 0 0
2
43232.7 0
0
7 74LS190
134 377 315 0 14 29
0 2 29 27 11 20 19 18 17 37
31 8 3 28 7
0
0 0 4336 0
7 74LS190
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
3656 0 0
2
43232.7 0
0
59
0 2 3 0 0 4096 0 0 6 52 0 4
537 487
537 512
540 512
540 525
1 6 4 0 0 4224 0 2 5 0 0 3
491 573
505 573
505 569
3 2 5 0 0 8320 0 3 2 0 0 3
457 571
457 573
473 573
2 3 6 0 0 4224 0 15 2 0 0 3
441 623
482 623
482 618
1 0 7 0 0 4096 0 3 0 0 50 2
466 519
466 502
2 0 8 0 0 4096 0 3 0 0 53 2
448 519
448 480
1 5 9 0 0 4224 0 4 5 0 0 3
528 532
528 535
526 535
2 0 2 0 0 4096 0 11 0 0 14 2
663 268
617 268
4 0 2 0 0 0 0 11 0 0 14 2
663 286
617 286
3 0 2 0 0 0 0 11 0 0 14 2
663 277
617 277
5 0 2 0 0 0 0 11 0 0 14 2
663 295
617 295
7 0 2 0 0 0 0 11 0 0 14 2
663 313
617 313
9 0 2 0 0 0 0 11 0 0 14 3
663 331
617 331
617 322
8 1 2 0 0 8320 0 11 8 0 0 3
663 322
617 322
617 213
1 6 10 0 0 4224 0 7 11 0 0 3
639 214
639 304
663 304
0 1 11 0 0 4096 0 0 11 45 0 3
484 234
663 234
663 259
1 10 2 0 0 0 0 9 11 0 0 3
652 349
652 340
657 340
1 10 2 0 0 0 0 10 14 0 0 3
312 537
312 521
314 521
2 0 2 0 0 0 0 14 0 0 30 2
320 449
250 449
4 0 2 0 0 0 0 14 0 0 30 3
320 467
250 467
250 458
6 0 12 0 0 4096 0 14 0 0 29 2
320 485
268 485
8 0 12 0 0 0 0 14 0 0 29 2
320 503
268 503
7 0 12 0 0 0 0 14 0 0 29 2
320 494
268 494
5 0 12 0 0 0 0 14 0 0 29 2
320 476
268 476
5 11 13 0 0 12416 0 19 11 0 0 6
525 330
513 330
513 384
742 384
742 277
727 277
12 6 14 0 0 12416 0 11 19 0 0 6
727 295
737 295
737 379
517 379
517 339
525 339
7 13 15 0 0 12416 0 19 11 0 0 6
525 348
521 348
521 375
732 375
732 313
727 313
8 14 16 0 0 8320 0 19 11 0 0 4
525 357
525 371
727 371
727 331
1 9 12 0 0 4224 0 12 14 0 0 3
268 443
268 512
320 512
3 1 2 0 0 0 0 14 13 0 0 3
320 458
250 458
250 441
1 0 11 0 0 0 0 14 0 0 45 3
320 440
278 440
278 315
14 8 17 0 0 8320 0 14 23 0 0 6
384 512
406 512
406 399
330 399
330 351
345 351
13 7 18 0 0 8320 0 14 23 0 0 6
384 494
398 494
398 407
323 407
323 342
345 342
12 6 19 0 0 16512 0 14 23 0 0 6
384 476
390 476
390 414
316 414
316 333
345 333
11 5 20 0 0 12416 0 14 23 0 0 5
384 458
384 420
310 420
310 324
345 324
1 0 21 0 0 4096 0 5 0 0 49 2
518 513
518 454
2 0 22 0 0 4096 0 5 0 0 48 2
509 513
509 460
3 0 23 0 0 4096 0 5 0 0 47 2
500 513
500 465
4 0 24 0 0 4096 0 5 0 0 46 2
491 513
491 472
1 3 25 0 0 8320 0 16 15 0 0 4
354 574
369 574
369 632
395 632
1 3 26 0 0 4224 0 15 6 0 0 3
441 641
549 641
549 570
0 3 27 0 0 4096 0 0 19 43 0 4
300 371
480 371
480 312
519 312
3 2 27 0 0 8320 0 23 16 0 0 4
339 306
300 306
300 574
318 574
0 1 22 0 0 4096 0 0 6 48 0 2
558 460
558 525
0 4 11 0 0 8320 0 0 19 58 0 5
278 315
278 234
485 234
485 321
525 321
4 11 24 0 0 12416 0 17 19 0 0 5
491 447
491 472
605 472
605 330
589 330
12 3 23 0 0 8320 0 19 17 0 0 5
589 339
600 339
600 465
497 465
497 447
13 2 22 0 0 8320 0 19 17 0 0 5
589 348
594 348
594 460
503 460
503 447
14 1 21 0 0 4224 0 19 17 0 0 4
589 357
589 454
509 454
509 447
14 1 7 0 0 8320 0 23 18 0 0 5
409 351
425 351
425 502
549 502
549 447
13 2 28 0 0 8320 0 23 18 0 0 5
409 342
431 342
431 494
543 494
543 447
12 3 3 0 0 8320 0 23 18 0 0 5
409 333
437 333
437 487
537 487
537 447
4 11 8 0 0 12416 0 18 23 0 0 5
531 447
531 480
444 480
444 324
409 324
0 2 29 0 0 8320 0 0 19 59 0 5
298 297
298 249
494 249
494 303
525 303
2 1 30 0 0 8320 0 20 19 0 0 3
477 315
477 294
519 294
10 1 31 0 0 4224 0 23 20 0 0 2
409 315
441 315
1 1 2 0 0 0 0 23 21 0 0 3
339 288
324 288
324 274
4 1 11 0 0 128 0 23 1 0 0 3
345 315
204 315
204 183
3 2 29 0 0 128 0 22 23 0 0 2
178 297
345 297
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
