CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
1013 88 1917 1018
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
1181 184 1294 281
42991634 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 593 818 0 1 11
0 35
0
0 0 21344 90
2 0V
11 0 25 8
5 Reset
8 -13 43 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89845e-315 0
0
13 Logic Switch~
5 653 55 0 1 11
0 32
0
0 0 21344 270
2 0V
-6 -22 8 -14
5 Clock
-16 -31 19 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89845e-315 0
0
13 Logic Switch~
5 167 337 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 x0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89845e-315 0
0
13 Logic Switch~
5 167 255 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 x1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89845e-315 0
0
14 Logic Display~
6 919 394 0 1 2
10 8
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 867 398 0 4 22
0 6 7 4 8
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 11 0
1 U
5572 0 0
2
5.89845e-315 0
0
8 4-In OR~
219 639 606 0 5 22
0 20 22 21 19 18
0
0 0 96 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 12 0
1 U
8901 0 0
2
5.89845e-315 0
0
8 4-In OR~
219 654 398 0 5 22
0 26 29 28 27 25
0
0 0 96 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
7361 0 0
2
5.89845e-315 0
0
9 4-In AND~
219 586 746 0 5 22
0 12 11 10 9 16
0
0 0 96 0
6 74LS21
-21 -28 21 -20
3 U8A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 10 0
1 U
4747 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 586 704 0 4 22
0 7 14 13 17
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 9 0
1 U
972 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 587 665 0 4 22
0 6 11 13 19
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 9 0
1 U
3472 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 587 627 0 4 22
0 6 11 14 21
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 9 0
1 U
9998 0 0
2
5.89845e-315 0
0
9 2-In AND~
219 587 589 0 3 22
0 12 7 22
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3536 0 0
2
5.89845e-315 0
0
9 2-In AND~
219 586 550 0 3 22
0 14 13 20
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4597 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 587 509 0 4 22
0 6 14 13 24
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 7 0
1 U
3835 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 586 457 0 4 22
0 30 10 9 27
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 7 0
1 U
3670 0 0
2
5.89845e-315 0
0
9 3-In AND~
219 589 291 0 4 22
0 5 10 9 33
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 7 0
1 U
5616 0 0
2
5.89845e-315 0
0
9 2-In AND~
219 587 421 0 3 22
0 12 5 28
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
9323 0 0
2
5.89845e-315 0
0
9 2-In AND~
219 586 384 0 3 22
0 12 10 29
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
317 0 0
2
5.89845e-315 0
0
9 2-In AND~
219 587 346 0 3 22
0 12 9 26
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3108 0 0
2
5.89845e-315 0
0
9 2-In AND~
219 589 248 0 3 22
0 7 5 34
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4299 0 0
2
5.89845e-315 0
0
8 2-In OR~
219 643 722 0 3 22
0 17 16 15
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
5.89845e-315 0
0
8 2-In OR~
219 652 491 0 3 22
0 5 24 23
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
7876 0 0
2
5.89845e-315 0
0
8 2-In OR~
219 653 260 0 3 22
0 34 33 31
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6369 0 0
2
5.89845e-315 0
0
7 Ground~
168 748 524 0 1 3
0 2
0
0 0 53344 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
5.89845e-315 0
0
7 Ground~
168 748 391 0 1 3
0 2
0
0 0 53344 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7100 0 0
2
5.89845e-315 0
0
7 Ground~
168 743 235 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
5.89845e-315 0
0
5 4027~
219 748 600 0 7 32
0 2 18 32 15 35 4 5
0
0 0 4704 0
4 4027
7 -60 35 -52
3 FF0
3 -60 24 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
7678 0 0
2
5.89845e-315 0
0
5 4027~
219 748 464 0 7 32
0 2 25 32 23 35 40 7
0
0 0 4704 0
4 4027
7 -60 35 -52
3 FF1
4 -61 25 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
961 0 0
2
5.89845e-315 0
0
5 4027~
219 743 307 0 7 32
0 2 31 32 7 35 41 6
0
0 0 4704 0
4 4027
7 -60 35 -52
3 FF2
3 -62 24 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3178 0 0
2
5.89845e-315 0
0
9 Inverter~
13 551 130 0 2 22
0 13 9
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3409 0 0
2
5.89845e-315 0
0
9 Inverter~
13 486 129 0 2 22
0 10 14
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3951 0 0
2
5.89845e-315 0
0
9 Inverter~
13 425 129 0 2 22
0 5 30
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
8885 0 0
2
5.89845e-315 0
0
9 Inverter~
13 363 128 0 2 22
0 7 11
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3780 0 0
2
5.89845e-315 0
0
9 Inverter~
13 301 128 0 2 22
0 6 12
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9265 0 0
2
5.89845e-315 0
0
84
0 0 3 0 0 8320 0 0 0 0 0 3
806 271
843 271
843 389
6 3 4 0 0 8320 0 28 6 0 0 3
778 582
843 582
843 407
7 0 5 0 0 8192 0 28 0 0 82 7
772 564
784 564
784 204
587 204
587 41
398 41
398 97
6 6 4 0 0 0 0 28 28 0 0 1
778 582
7 0 6 0 0 4096 0 30 0 0 7 2
767 271
771 271
0 0 7 0 0 16384 0 0 0 9 83 6
777 428
777 211
578 211
578 50
336 50
336 96
1 0 6 0 0 24576 0 6 0 0 84 8
843 389
843 271
771 271
771 220
570 220
570 61
274 61
274 96
1 4 8 0 0 4224 0 5 6 0 0 2
903 398
888 398
2 7 7 0 0 0 0 6 29 0 0 4
843 398
834 398
834 428
772 428
4 0 9 0 0 4096 0 9 0 0 71 2
562 760
554 760
3 0 10 0 0 4096 0 9 0 0 81 2
562 751
459 751
2 0 11 0 0 4096 0 9 0 0 68 2
562 742
366 742
1 0 12 0 0 4096 0 9 0 0 67 2
562 733
304 733
3 0 13 0 0 4096 0 10 0 0 80 2
562 713
528 713
2 0 14 0 0 4096 0 10 0 0 70 2
562 704
489 704
1 0 7 0 0 0 0 10 0 0 83 2
562 695
336 695
3 4 15 0 0 8320 0 22 28 0 0 4
676 722
695 722
695 582
724 582
5 2 16 0 0 8320 0 9 22 0 0 4
607 746
618 746
618 731
630 731
4 1 17 0 0 12416 0 10 22 0 0 4
607 704
617 704
617 713
630 713
3 0 13 0 0 4096 0 11 0 0 80 2
563 674
528 674
2 0 11 0 0 4096 0 11 0 0 68 2
563 665
366 665
1 0 6 0 0 0 0 11 0 0 84 2
563 656
274 656
3 0 14 0 0 4096 0 12 0 0 70 2
563 636
489 636
2 0 11 0 0 0 0 12 0 0 68 2
563 627
366 627
1 0 6 0 0 0 0 12 0 0 84 2
563 618
274 618
2 0 7 0 0 0 0 13 0 0 83 2
563 598
336 598
1 0 12 0 0 4096 0 13 0 0 67 2
563 580
304 580
2 0 13 0 0 0 0 14 0 0 80 2
562 559
528 559
1 0 14 0 0 0 0 14 0 0 70 2
562 541
489 541
5 2 18 0 0 8320 0 7 28 0 0 4
672 606
682 606
682 564
724 564
4 4 19 0 0 8320 0 11 7 0 0 4
608 665
616 665
616 620
622 620
3 1 20 0 0 8320 0 14 7 0 0 4
607 550
616 550
616 593
622 593
4 3 21 0 0 4224 0 12 7 0 0 3
608 627
608 611
622 611
3 2 22 0 0 8320 0 13 7 0 0 3
608 589
608 602
622 602
3 0 13 0 0 0 0 15 0 0 80 2
563 518
528 518
2 0 14 0 0 0 0 15 0 0 70 2
563 509
489 509
1 0 6 0 0 0 0 15 0 0 84 2
563 500
274 500
3 4 23 0 0 4224 0 23 29 0 0 3
685 491
685 446
724 446
4 2 24 0 0 12416 0 15 23 0 0 4
608 509
616 509
616 500
639 500
1 0 5 0 0 0 0 23 0 0 82 2
639 482
398 482
5 2 25 0 0 8320 0 8 29 0 0 4
687 398
694 398
694 428
724 428
3 1 26 0 0 8320 0 20 8 0 0 4
608 346
626 346
626 385
637 385
4 4 27 0 0 8320 0 16 8 0 0 4
607 457
624 457
624 412
637 412
3 3 28 0 0 12416 0 18 8 0 0 4
608 421
614 421
614 403
637 403
3 2 29 0 0 12416 0 19 8 0 0 4
607 384
613 384
613 394
637 394
3 0 9 0 0 0 0 16 0 0 71 2
562 466
554 466
2 0 10 0 0 0 0 16 0 0 81 2
562 457
459 457
1 0 30 0 0 4096 0 16 0 0 69 2
562 448
428 448
2 0 5 0 0 0 0 18 0 0 82 2
563 430
398 430
1 0 12 0 0 0 0 18 0 0 67 2
563 412
304 412
2 0 10 0 0 0 0 19 0 0 81 2
562 393
459 393
1 0 12 0 0 0 0 19 0 0 67 2
562 375
304 375
2 0 9 0 0 4096 0 20 0 0 71 2
563 355
554 355
1 0 12 0 0 0 0 20 0 0 67 2
563 337
304 337
4 0 7 0 0 12288 0 30 0 0 83 4
719 289
655 289
655 317
336 317
3 2 31 0 0 8320 0 24 30 0 0 3
686 260
686 271
719 271
3 0 32 0 0 4096 0 30 0 0 59 2
719 280
706 280
3 0 32 0 0 4096 0 29 0 0 59 2
724 437
706 437
1 3 32 0 0 12416 0 2 28 0 0 5
653 67
653 128
706 128
706 573
724 573
4 2 33 0 0 4224 0 17 24 0 0 4
610 291
632 291
632 269
640 269
3 1 34 0 0 4224 0 21 24 0 0 4
610 248
632 248
632 251
640 251
3 0 9 0 0 4096 0 17 0 0 71 2
565 300
554 300
2 0 10 0 0 4096 0 17 0 0 81 2
565 291
459 291
1 0 5 0 0 0 0 17 0 0 82 2
565 282
398 282
2 0 5 0 0 0 0 21 0 0 82 2
565 257
398 257
1 0 7 0 0 0 0 21 0 0 83 2
565 239
336 239
2 0 12 0 0 4224 0 35 0 0 0 2
304 146
304 772
2 0 11 0 0 4224 0 34 0 0 0 2
366 146
366 772
2 0 30 0 0 4224 0 33 0 0 0 2
428 147
428 772
2 0 14 0 0 4224 0 32 0 0 0 2
489 147
489 774
2 0 9 0 0 4224 0 31 0 0 0 2
554 148
554 775
5 0 35 0 0 8192 0 28 0 0 74 3
748 606
748 636
716 636
5 0 35 0 0 0 0 29 0 0 74 3
748 470
748 493
716 493
1 5 35 0 0 12416 0 1 30 0 0 6
594 805
594 776
716 776
716 329
743 329
743 313
1 1 2 0 0 4224 0 28 25 0 0 2
748 543
748 532
1 1 2 0 0 0 0 26 29 0 0 2
748 399
748 407
1 1 2 0 0 0 0 27 30 0 0 2
743 243
743 250
1 0 10 0 0 12288 0 4 0 0 81 5
179 255
242 255
242 71
459 71
459 98
1 0 13 0 0 12288 0 3 0 0 80 5
179 337
253 337
253 82
528 82
528 100
1 0 13 0 0 12416 0 31 0 0 0 4
554 112
554 100
528 100
528 774
1 0 10 0 0 12416 0 32 0 0 0 4
489 111
489 98
459 98
459 774
1 0 5 0 0 12416 0 33 0 0 0 4
428 111
428 97
398 97
398 773
1 0 7 0 0 12416 0 34 0 0 0 4
366 110
366 96
336 96
336 772
1 0 6 0 0 12416 0 35 0 0 0 4
304 110
304 96
274 96
274 773
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
