CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 100 10
775 149 1679 1079
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
943 245 1056 342
42991634 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 685 180 0 1 11
0 18
0
0 0 21360 270
2 0V
-6 -21 8 -13
5 Reset
-16 -31 19 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89846e-315 0
0
13 Logic Switch~
5 99 116 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 Modo
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89846e-315 0
0
9 Inverter~
13 194 411 0 2 22
0 3 6
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U4E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3124 0 0
2
5.89846e-315 0
0
9 2-In AND~
219 189 352 0 3 22
0 4 6 5
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U9A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3421 0 0
2
5.89846e-315 0
0
5 4073~
219 303 437 0 4 22
0 9 10 8 7
0
0 0 624 270
4 4073
-7 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
8157 0 0
2
5.89846e-315 0
0
9 2-In AND~
219 303 363 0 3 22
0 11 12 10
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5572 0 0
2
5.89846e-315 0
0
5 4025~
219 354 353 0 4 22
0 13 14 15 9
0
0 0 624 270
4 4025
-14 -24 14 -16
3 U7A
31 -10 52 -2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 5 0
1 U
8901 0 0
2
5.89846e-315 0
0
8 2-In OR~
219 119 318 0 3 22
0 5 16 4
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U8A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7361 0 0
2
5.89846e-315 0
0
8 3-In OR~
219 641 268 0 4 22
0 7 17 18 3
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U6A
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
4747 0 0
2
5.89846e-315 0
0
9 Inverter~
13 404 312 0 2 22
0 8 19
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U4D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
972 0 0
2
5.89846e-315 0
0
5 4073~
219 439 357 0 4 22
0 13 15 19 17
0
0 0 624 270
4 4073
-7 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
3472 0 0
2
5.89846e-315 0
0
2 +V
167 255 247 0 1 3
0 20
0
0 0 53488 90
2 5V
-7 -15 7 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.89846e-315 0
0
7 Ground~
168 256 224 0 1 3
0 2
0
0 0 53360 270
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.89846e-315 0
0
7 Ground~
168 490 227 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89846e-315 0
0
12 Hex Display~
7 419 115 0 16 19
10 13 23 22 21 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3835 0 0
2
5.89846e-315 0
0
12 Hex Display~
7 457 115 0 18 19
10 14 11 12 15 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3670 0 0
2
5.89846e-315 0
0
9 2-In AND~
219 173 171 0 3 22
0 8 16 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5616 0 0
2
5.89846e-315 0
0
9 Inverter~
13 224 171 0 2 22
0 28 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9323 0 0
2
5.89846e-315 0
0
9 Inverter~
13 263 153 0 2 22
0 26 25
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
317 0 0
2
5.89846e-315 0
0
9 Inverter~
13 178 116 0 2 22
0 8 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3108 0 0
2
5.89846e-315 0
0
9 2-In AND~
219 239 125 0 3 22
0 27 16 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4299 0 0
2
5.89846e-315 0
0
7 Pulser~
4 65 189 0 10 12
0 31 32 16 33 0 0 10 10 10
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9672 0 0
2
5.89846e-315 0
0
7 74LS193
137 546 210 0 14 29
0 30 29 5 3 2 2 2 8 34
35 21 22 23 13
0
0 0 4336 0
7 74LS193
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
5.89846e-315 0
0
7 74LS193
137 312 209 0 14 29
0 25 24 5 3 2 20 20 20 30
29 15 12 11 14
0
0 0 4336 0
7 74LS193
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
5.89846e-315 0
0
51
1 0 3 0 0 8192 0 3 0 0 23 3
197 429
251 429
251 268
1 3 4 0 0 4224 0 4 8 0 0 3
179 373
122 373
122 348
1 0 5 0 0 8192 0 8 0 0 4 3
131 302
131 289
188 289
3 0 5 0 0 4096 0 4 0 0 24 3
188 328
188 227
200 227
2 2 6 0 0 4224 0 4 3 0 0 2
197 373
197 393
4 1 7 0 0 4224 0 5 9 0 0 4
301 460
674 460
674 277
660 277
3 0 8 0 0 12288 0 5 0 0 32 4
292 415
292 390
264 390
264 278
1 4 9 0 0 8320 0 5 7 0 0 4
310 415
310 390
360 390
360 386
3 2 10 0 0 4224 0 6 5 0 0 2
301 386
301 415
1 0 11 0 0 8192 0 6 0 0 39 4
310 341
310 313
388 313
388 236
2 0 12 0 0 8192 0 6 0 0 38 4
292 341
292 304
378 304
378 227
1 0 13 0 0 8192 0 7 0 0 18 3
369 334
369 286
446 286
2 0 14 0 0 4096 0 7 0 0 40 2
360 335
360 245
3 0 15 0 0 4096 0 7 0 0 37 2
351 334
351 218
0 2 16 0 0 4224 0 0 8 41 0 2
113 180
113 302
2 4 17 0 0 12416 0 9 11 0 0 4
659 268
685 268
685 380
437 380
3 1 18 0 0 8320 0 9 1 0 0 3
660 259
685 259
685 192
1 0 13 0 0 8192 0 11 0 0 36 4
446 335
446 286
587 286
587 246
2 0 15 0 0 4224 0 11 0 0 37 2
437 335
437 218
2 3 19 0 0 8320 0 10 11 0 0 3
407 330
407 335
428 335
1 0 8 0 0 0 0 10 0 0 32 2
407 294
407 278
0 4 3 0 0 0 0 0 9 23 0 2
477 268
614 268
4 4 3 0 0 12416 0 24 23 0 0 6
280 209
239 209
239 268
477 268
477 210
514 210
3 3 5 0 0 12416 0 23 24 0 0 6
508 201
472 201
472 259
200 259
200 200
274 200
7 0 20 0 0 4096 0 24 0 0 26 2
280 236
272 236
6 0 20 0 0 8320 0 24 0 0 27 3
280 227
272 227
272 245
1 8 20 0 0 0 0 12 24 0 0 2
266 245
280 245
1 5 2 0 0 12288 0 13 24 0 0 4
263 225
268 225
268 218
280 218
5 0 2 0 0 0 0 23 0 0 30 3
514 219
506 219
506 229
7 0 2 0 0 0 0 23 0 0 31 3
514 237
506 237
506 228
1 6 2 0 0 4224 0 14 23 0 0 2
497 228
514 228
8 0 8 0 0 12416 0 23 0 0 48 5
514 246
497 246
497 278
129 278
129 160
11 4 21 0 0 12416 0 23 15 0 0 5
578 219
603 219
603 162
410 162
410 139
12 3 22 0 0 12416 0 23 15 0 0 5
578 228
598 228
598 157
416 157
416 139
13 2 23 0 0 12416 0 23 15 0 0 5
578 237
593 237
593 152
422 152
422 139
14 1 13 0 0 12416 0 23 15 0 0 5
578 246
588 246
588 147
428 147
428 139
11 4 15 0 0 0 0 24 16 0 0 3
344 218
448 218
448 139
12 3 12 0 0 4224 0 24 16 0 0 3
344 227
454 227
454 139
13 2 11 0 0 4224 0 24 16 0 0 3
344 236
460 236
460 139
1 14 14 0 0 8320 0 16 24 0 0 3
466 139
466 245
344 245
2 0 16 0 0 0 0 21 0 0 42 3
215 134
113 134
113 180
3 2 16 0 0 0 0 22 17 0 0 2
89 180
149 180
2 2 24 0 0 12416 0 18 24 0 0 4
245 171
254 171
254 191
280 191
2 1 25 0 0 8320 0 19 24 0 0 3
266 171
266 182
280 182
3 1 26 0 0 8320 0 21 19 0 0 3
260 125
266 125
266 135
2 1 27 0 0 4224 0 20 21 0 0 2
199 116
215 116
1 0 8 0 0 0 0 20 0 0 48 2
163 116
129 116
1 1 8 0 0 0 0 2 17 0 0 4
111 116
129 116
129 162
149 162
3 1 28 0 0 4224 0 17 18 0 0 2
194 171
209 171
10 2 29 0 0 4224 0 24 23 0 0 4
350 209
439 209
439 192
514 192
9 1 30 0 0 12416 0 24 23 0 0 4
350 200
430 200
430 183
514 183
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
