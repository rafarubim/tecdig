CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
1180 88 1917 1018
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
1348 184 1461 281
42991634 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 519 582 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
6 Ligado
-3 -10 39 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9730 0 0
2
43178.2 0
0
13 Logic Switch~
5 268 629 0 1 11
0 12
0
0 0 21360 90
2 0V
11 0 25 8
1 E
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9874 0 0
2
5.89839e-315 0
0
13 Logic Switch~
5 214 628 0 1 11
0 13
0
0 0 21360 90
2 0V
11 0 25 8
1 D
13 -10 20 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
364 0 0
2
5.89839e-315 0
0
13 Logic Switch~
5 159 627 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
1 C
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3656 0 0
2
5.89839e-315 0
0
13 Logic Switch~
5 106 626 0 1 11
0 15
0
0 0 21360 90
2 0V
11 0 25 8
1 B
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3131 0 0
2
5.89839e-315 0
0
13 Logic Switch~
5 60 624 0 1 11
0 16
0
0 0 21360 90
2 0V
11 0 25 8
1 A
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6772 0 0
2
5.89839e-315 0
0
5 4068~
219 544 416 0 9 19
0 10 9 8 7 6 5 4 3 11
0
0 0 624 0
4 4068
-7 -24 21 -16
2 U3
-8 -44 6 -36
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 0 0 0 0
1 U
9557 0 0
2
43178.2 0
0
5 4023~
219 400 543 0 4 22
0 16 15 13 4
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 9 0
1 U
5789 0 0
2
43178.2 0
0
5 4023~
219 401 496 0 4 22
0 16 15 14 5
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 9 0
1 U
7328 0 0
2
43178.2 0
0
5 4023~
219 400 396 0 4 22
0 15 19 13 7
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 9 0
1 U
4799 0 0
2
43178.2 0
0
10 4-In NAND~
219 401 449 0 5 22
0 16 20 19 12 6
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U1B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 8 0
1 U
9196 0 0
2
43178.2 0
0
10 4-In NAND~
219 401 341 0 5 22
0 21 19 13 17 8
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U1A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 8 0
1 U
3857 0 0
2
43178.2 0
0
10 4-In NAND~
219 400 288 0 5 22
0 21 15 18 12 9
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U7B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
7125 0 0
2
43178.2 0
0
10 4-In NAND~
219 400 236 0 5 22
0 21 20 19 18 10
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U7A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
3641 0 0
2
43178.2 0
0
5 4049~
219 255 453 0 2 22
0 12 17
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4E
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
9821 0 0
2
5.89839e-315 0
0
5 4049~
219 200 481 0 2 22
0 13 18
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4D
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
3187 0 0
2
5.89839e-315 0
0
5 4049~
219 147 443 0 2 22
0 14 19
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4C
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
762 0 0
2
5.89839e-315 0
0
5 4049~
219 95 482 0 2 22
0 15 20
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4B
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
39 0 0
2
5.89839e-315 0
0
5 4049~
219 60 438 0 2 22
0 16 21
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4A
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
9450 0 0
2
5.89839e-315 0
0
7 Ground~
168 619 416 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3236 0 0
2
5.89839e-315 0
0
4 LED~
171 587 415 0 2 2
10 11 2
0
0 0 864 90
4 LED1
-12 -21 16 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3321 0 0
2
5.89839e-315 0
0
42
8 1 3 0 0 4224 0 7 1 0 0 2
520 448
520 569
4 7 4 0 0 8320 0 8 7 0 0 4
427 543
502 543
502 439
520 439
4 6 5 0 0 4224 0 9 7 0 0 4
428 496
507 496
507 430
520 430
5 5 6 0 0 4224 0 11 7 0 0 4
428 449
512 449
512 421
520 421
4 4 7 0 0 4224 0 10 7 0 0 4
427 396
512 396
512 412
520 412
5 3 8 0 0 4224 0 12 7 0 0 4
428 341
502 341
502 403
520 403
5 2 9 0 0 8320 0 13 7 0 0 4
427 288
507 288
507 394
520 394
5 1 10 0 0 8320 0 14 7 0 0 4
427 236
512 236
512 385
520 385
2 1 2 0 0 8320 0 21 20 0 0 3
600 416
600 417
612 417
9 1 11 0 0 8320 0 7 21 0 0 3
571 416
571 416
580 416
4 0 12 0 0 4096 0 11 0 0 12 2
377 463
325 463
0 4 12 0 0 16512 0 0 13 38 0 6
258 571
269 571
269 572
325 572
325 302
376 302
3 0 13 0 0 4096 0 8 0 0 15 3
376 552
280 552
280 535
3 0 13 0 0 0 0 10 0 0 15 2
376 405
280 405
0 3 13 0 0 12416 0 0 12 39 0 5
203 536
203 535
280 535
280 346
377 346
0 0 14 0 0 8192 0 0 0 17 40 3
165 524
165 525
151 525
0 3 14 0 0 4224 0 0 9 0 0 4
159 524
313 524
313 505
377 505
2 0 15 0 0 4096 0 8 0 0 22 5
376 543
315 543
315 542
305 542
305 514
0 2 15 0 0 4096 0 0 9 22 0 4
305 497
370 497
370 496
377 496
0 1 15 0 0 4096 0 0 10 22 0 2
305 387
376 387
0 0 15 0 0 0 0 0 0 22 41 3
106 514
106 515
98 515
0 2 15 0 0 8320 0 0 13 0 0 4
103 514
305 514
305 284
376 284
1 0 16 0 0 4096 0 8 0 0 25 3
376 534
298 534
298 506
1 0 16 0 0 4096 0 9 0 0 25 2
377 487
298 487
0 1 16 0 0 4224 0 0 11 42 0 4
63 506
298 506
298 436
377 436
2 4 17 0 0 16512 0 15 12 0 0 5
258 435
258 427
259 427
259 355
377 355
3 0 18 0 0 4096 0 13 0 0 28 4
376 293
208 293
208 294
203 294
2 4 18 0 0 4224 0 16 14 0 0 3
203 463
203 250
376 250
3 0 19 0 0 16384 0 11 0 0 30 5
377 454
372 454
372 453
333 453
333 396
2 0 19 0 0 4224 0 10 0 0 32 2
376 396
151 396
2 0 19 0 0 4224 0 12 0 0 32 2
377 337
151 337
2 3 19 0 0 0 0 17 14 0 0 4
150 425
151 425
151 241
376 241
2 0 20 0 0 20480 0 11 0 0 34 6
377 445
368 445
368 446
292 446
292 412
98 412
2 2 20 0 0 8320 0 18 14 0 0 3
98 464
98 232
376 232
1 0 21 0 0 4224 0 12 0 0 37 2
377 328
62 328
1 0 21 0 0 0 0 13 0 0 37 2
376 275
62 275
2 1 21 0 0 0 0 19 14 0 0 5
63 420
63 390
62 390
62 223
376 223
1 1 12 0 0 0 0 15 2 0 0 4
258 471
258 609
269 609
269 616
1 1 13 0 0 0 0 16 3 0 0 4
203 499
203 608
215 608
215 615
1 1 14 0 0 0 0 17 4 0 0 5
150 461
151 461
151 607
160 607
160 614
1 1 15 0 0 0 0 18 5 0 0 4
98 500
98 606
107 606
107 613
1 1 16 0 0 0 0 19 6 0 0 4
63 456
63 604
61 604
61 611
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
