CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 21 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
8
9 2-In AND~
219 676 459 0 3 22
0 5 4 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9172 0 0
2
43198.6 0
0
12 Hex Display~
7 594 521 0 18 19
10 5 4 11 10 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7100 0 0
2
43198.6 0
0
12 Hex Display~
7 552 521 0 16 19
10 9 6 8 7 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3820 0 0
2
43198.6 1
0
7 Ground~
168 697 322 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
43198.6 3
0
7 74LS290
153 729 384 0 10 21
0 2 2 3 6 8 10 8 6 9
7
0
0 0 4336 0
7 74LS290
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
961 0 0
2
43198.6 4
0
7 Ground~
168 561 320 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
43198.6 5
0
7 74LS290
153 593 384 0 10 21
0 2 2 3 6 11 12 11 4 5
10
0
0 0 4336 0
7 74LS290
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
3409 0 0
2
43198.6 6
0
7 Pulser~
4 467 420 0 10 12
0 13 14 12 15 0 0 30 30 17
7
0
0 0 4144 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3951 0 0
2
43198.6 7
0
22
0 3 3 0 0 4224 0 0 7 2 0 4
680 435
545 435
545 375
561 375
3 3 3 0 0 0 0 1 5 0 0 5
697 459
697 435
679 435
679 375
697 375
2 0 4 0 0 4096 0 1 0 0 13 2
652 468
637 468
1 0 5 0 0 4096 0 1 0 0 14 2
652 450
632 450
0 4 6 0 0 4096 0 0 7 6 0 4
685 425
550 425
550 384
561 384
0 4 6 0 0 0 0 0 5 9 0 4
774 425
685 425
685 384
697 384
10 4 7 0 0 8320 0 5 3 0 0 4
761 411
761 589
543 589
543 545
7 3 8 0 0 12416 0 5 3 0 0 5
761 357
780 357
780 583
549 583
549 545
8 2 6 0 0 12416 0 5 3 0 0 5
761 375
774 375
774 576
555 576
555 545
9 1 9 0 0 12416 0 5 3 0 0 5
761 393
768 393
768 569
561 569
561 545
4 0 10 0 0 12416 0 2 0 0 17 4
585 545
585 563
647 563
647 411
7 3 11 0 0 8320 0 7 2 0 0 5
625 357
642 357
642 557
591 557
591 545
8 2 4 0 0 8320 0 7 2 0 0 5
625 375
637 375
637 552
597 552
597 545
9 1 5 0 0 8320 0 7 2 0 0 4
625 393
632 393
632 545
603 545
7 5 8 0 0 0 0 5 5 0 0 5
761 357
761 306
669 306
669 402
691 402
5 7 11 0 0 0 0 7 7 0 0 5
555 402
539 402
539 306
625 306
625 357
10 6 10 0 0 0 0 7 5 0 0 2
625 411
691 411
3 6 12 0 0 4224 0 8 7 0 0 2
491 411
555 411
1 1 2 0 0 4096 0 5 4 0 0 2
697 357
697 330
2 1 2 0 0 0 0 5 5 0 0 2
697 366
697 357
1 1 2 0 0 4224 0 7 6 0 0 2
561 357
561 328
2 1 2 0 0 0 0 7 7 0 0 2
561 366
561 357
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
