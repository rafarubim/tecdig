CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 42 379 0 1 11
0 42
0
0 0 21360 90
2 0V
11 0 25 8
1 E
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4484 0 0
2
5.89841e-315 0
0
13 Logic Switch~
5 217 623 0 1 11
0 38
0
0 0 21360 90
2 0V
11 0 25 8
2 C0
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5996 0 0
2
5.89841e-315 0
0
13 Logic Switch~
5 177 622 0 1 11
0 39
0
0 0 21360 90
2 0V
11 0 25 8
2 C1
12 -10 26 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7804 0 0
2
5.89841e-315 0
0
13 Logic Switch~
5 138 621 0 1 11
0 40
0
0 0 21360 90
2 0V
11 0 25 8
2 C2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5523 0 0
2
5.89841e-315 0
0
13 Logic Switch~
5 99 620 0 1 11
0 41
0
0 0 21360 90
2 0V
11 0 25 8
2 C3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3330 0 0
2
5.89841e-315 0
0
9 Inverter~
13 421 619 0 2 22
0 18 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3465 0 0
2
43192 0
0
9 Inverter~
13 416 574 0 2 22
0 19 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
8396 0 0
2
43192 0
0
9 Inverter~
13 420 540 0 2 22
0 20 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3685 0 0
2
43192 0
0
9 Inverter~
13 416 499 0 2 22
0 21 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
7849 0 0
2
43192 0
0
9 Inverter~
13 416 461 0 2 22
0 22 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
6343 0 0
2
43192 0
0
9 Inverter~
13 423 424 0 2 22
0 23 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
7376 0 0
2
43192 0
0
9 Inverter~
13 429 388 0 2 22
0 24 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
9156 0 0
2
43192 0
0
9 Inverter~
13 435 351 0 2 22
0 25 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
5776 0 0
2
43192 0
0
9 Inverter~
13 425 312 0 2 22
0 26 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
7207 0 0
2
43192 0
0
9 Inverter~
13 428 273 0 2 22
0 27 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4459 0 0
2
43192 0
0
9 Inverter~
13 433 238 0 2 22
0 28 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3760 0 0
2
43192 0
0
9 Inverter~
13 440 207 0 2 22
0 29 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
754 0 0
2
43192 0
0
9 Inverter~
13 443 156 0 2 22
0 30 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9767 0 0
2
43192 0
0
9 Inverter~
13 449 122 0 2 22
0 31 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
7978 0 0
2
43192 0
0
9 Inverter~
13 448 88 0 2 22
0 32 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3142 0 0
2
43192 0
0
9 Inverter~
13 446 50 0 2 22
0 33 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3284 0 0
2
43192 0
0
14 Logic Display~
6 473 616 0 1 2
10 2
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L16
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
659 0 0
2
5.89841e-315 5.42414e-315
0
14 Logic Display~
6 470 570 0 1 2
10 3
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L15
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
5.89841e-315 5.41896e-315
0
14 Logic Display~
6 472 536 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L14
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6792 0 0
2
5.89841e-315 5.41378e-315
0
14 Logic Display~
6 477 495 0 1 2
10 5
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L13
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
5.89841e-315 5.4086e-315
0
14 Logic Display~
6 476 456 0 1 2
10 6
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L12
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6316 0 0
2
5.89841e-315 5.40342e-315
0
14 Logic Display~
6 478 421 0 1 2
10 7
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L11
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8734 0 0
2
5.89841e-315 5.39824e-315
0
14 Logic Display~
6 483 384 0 1 2
10 8
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L10
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7988 0 0
2
5.89841e-315 5.39306e-315
0
14 Logic Display~
6 488 348 0 1 2
10 9
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L9
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3217 0 0
2
5.89841e-315 5.38788e-315
0
14 Logic Display~
6 487 308 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3965 0 0
2
5.89841e-315 5.37752e-315
0
14 Logic Display~
6 488 269 0 1 2
10 11
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8239 0 0
2
5.89841e-315 5.36716e-315
0
14 Logic Display~
6 493 235 0 1 2
10 12
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
828 0 0
2
5.89841e-315 5.3568e-315
0
14 Logic Display~
6 498 203 0 1 2
10 13
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
5.89841e-315 5.34643e-315
0
14 Logic Display~
6 496 152 0 1 2
10 14
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7107 0 0
2
5.89841e-315 5.32571e-315
0
14 Logic Display~
6 499 111 0 1 2
10 15
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6433 0 0
2
5.89841e-315 5.30499e-315
0
14 Logic Display~
6 500 84 0 1 2
10 16
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8559 0 0
2
5.89841e-315 5.26354e-315
0
14 Logic Display~
6 499 58 0 1 2
10 17
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3674 0 0
2
5.89841e-315 0
0
7 74LS139
118 330 547 0 14 29
0 39 38 34 43 44 45 21 20 19
18 46 47 48 49
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
5697 0 0
2
5.89841e-315 0
0
7 74LS139
118 328 401 0 14 29
0 39 38 35 50 51 52 25 24 23
22 53 54 55 56
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
3805 0 0
2
5.89841e-315 0
0
7 74LS139
118 326 248 0 14 29
0 39 38 36 57 58 59 29 28 27
26 60 61 62 63
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
5219 0 0
2
5.89841e-315 0
0
7 74LS139
118 325 89 0 14 29
0 39 38 37 64 65 66 33 32 31
30 67 68 69 70
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
3795 0 0
2
5.89841e-315 0
0
7 74LS139
118 149 315 0 14 29
0 41 40 42 71 72 73 37 36 35
34 74 75 76 77
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
3637 0 0
2
5.89841e-315 0
0
47
2 1 2 0 0 8320 0 6 22 0 0 3
442 619
442 620
457 620
2 1 3 0 0 4224 0 7 23 0 0 2
437 574
454 574
2 1 4 0 0 4224 0 8 24 0 0 2
441 540
456 540
2 1 5 0 0 4224 0 9 25 0 0 2
437 499
461 499
2 1 6 0 0 8320 0 10 26 0 0 3
437 461
437 460
460 460
2 1 7 0 0 8320 0 11 27 0 0 3
444 424
444 425
462 425
2 1 8 0 0 4224 0 12 28 0 0 2
450 388
467 388
2 1 9 0 0 8320 0 13 29 0 0 3
456 351
456 352
472 352
2 1 10 0 0 4224 0 14 30 0 0 2
446 312
471 312
2 1 11 0 0 4224 0 15 31 0 0 2
449 273
472 273
2 1 12 0 0 8320 0 16 32 0 0 3
454 238
454 239
477 239
2 1 13 0 0 4224 0 17 33 0 0 2
461 207
482 207
2 1 14 0 0 4224 0 18 34 0 0 2
464 156
480 156
2 1 15 0 0 8320 0 19 35 0 0 4
470 122
476 122
476 115
483 115
2 1 16 0 0 4224 0 20 36 0 0 2
469 88
484 88
2 1 17 0 0 8320 0 21 37 0 0 4
467 50
474 50
474 62
483 62
10 1 18 0 0 8320 0 38 6 0 0 5
368 547
377 547
377 620
406 620
406 619
9 1 19 0 0 8320 0 38 7 0 0 4
368 538
383 538
383 574
401 574
8 1 20 0 0 4224 0 38 8 0 0 4
368 529
389 529
389 540
405 540
7 1 21 0 0 8320 0 38 9 0 0 4
368 520
383 520
383 499
401 499
10 1 22 0 0 8320 0 39 10 0 0 5
366 401
371 401
371 460
401 460
401 461
9 1 23 0 0 8320 0 39 11 0 0 5
366 392
378 392
378 425
408 425
408 424
8 1 24 0 0 12416 0 39 12 0 0 4
366 383
386 383
386 388
414 388
7 1 25 0 0 12416 0 39 13 0 0 5
366 374
386 374
386 352
420 352
420 351
10 1 26 0 0 8320 0 40 14 0 0 4
364 248
369 248
369 312
410 312
9 1 27 0 0 12416 0 40 15 0 0 4
364 239
377 239
377 273
413 273
8 1 28 0 0 12416 0 40 16 0 0 5
364 230
385 230
385 239
418 239
418 238
7 1 29 0 0 12416 0 40 17 0 0 4
364 221
377 221
377 207
425 207
10 1 30 0 0 8320 0 41 18 0 0 4
363 89
371 89
371 156
428 156
9 1 31 0 0 12416 0 41 19 0 0 4
363 80
381 80
381 122
434 122
8 1 32 0 0 12416 0 41 20 0 0 4
363 71
390 71
390 88
433 88
7 1 33 0 0 12416 0 41 21 0 0 4
363 62
378 62
378 50
431 50
10 3 34 0 0 8320 0 42 38 0 0 4
187 315
244 315
244 547
292 547
9 3 35 0 0 8320 0 42 39 0 0 4
187 306
267 306
267 401
290 401
8 3 36 0 0 4224 0 42 40 0 0 4
187 297
267 297
267 248
288 248
7 3 37 0 0 8320 0 42 41 0 0 4
187 288
244 288
244 89
287 89
2 0 38 0 0 4096 0 40 0 0 44 2
294 239
218 239
2 0 38 0 0 4096 0 39 0 0 44 2
296 392
218 392
2 0 38 0 0 4096 0 38 0 0 44 2
298 538
218 538
1 0 39 0 0 4096 0 40 0 0 43 2
294 230
213 230
1 0 39 0 0 4096 0 39 0 0 43 2
296 383
213 383
1 0 39 0 0 4096 0 38 0 0 43 2
298 529
213 529
1 1 39 0 0 12416 0 3 41 0 0 5
178 609
178 587
213 587
213 71
293 71
1 2 38 0 0 4224 0 2 41 0 0 3
218 610
218 80
293 80
1 2 40 0 0 12416 0 4 42 0 0 5
139 608
139 587
105 587
105 306
117 306
1 1 41 0 0 4224 0 5 42 0 0 3
100 607
100 297
117 297
1 3 42 0 0 8320 0 1 42 0 0 3
43 366
43 315
111 315
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
