CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
238 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
406 176 519 273
42991634 0
0
6 Title:
5 Name:
0
0
0
47
13 Logic Switch~
5 773 443 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
5 Reset
-16 -31 19 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7376 0 0
2
43239.8 0
0
9 Inverter~
13 689 562 0 2 22
0 4 3
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U12D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
9156 0 0
2
43239.8 0
0
9 Inverter~
13 645 562 0 2 22
0 5 4
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U12C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
5776 0 0
2
43239.8 0
0
9 Inverter~
13 602 562 0 2 22
0 6 5
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U12B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
7207 0 0
2
43239.8 0
0
9 Inverter~
13 555 562 0 2 22
0 8 6
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U12A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
4459 0 0
2
43239.8 0
0
12 Hex Display~
7 897 485 0 16 19
10 12 11 10 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3760 0 0
2
43239.8 0
0
7 74LS175
131 817 568 0 14 29
0 7 3 13 14 15 16 9 47 10
48 11 49 12 50
0
0 0 4336 0
7 74LS175
-24 -51 25 -43
3 U11
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
754 0 0
2
43239.8 0
0
8 2-In OR~
219 162 750 0 3 22
0 18 8 17
0
0 0 112 90
6 74LS32
-21 -24 21 -16
4 U10A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9767 0 0
2
43239.8 0
0
9 2-In AND~
219 698 708 0 3 22
0 20 22 16
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U7B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7978 0 0
2
43239.8 4
0
9 2-In AND~
219 698 672 0 3 22
0 20 19 15
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U7A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3142 0 0
2
43239.8 3
0
10 3-In NAND~
219 589 644 0 4 22
0 22 19 21 20
0
0 0 112 90
6 74LS10
-21 -28 21 -20
3 U8A
19 -2 40 6
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
3284 0 0
2
43239.8 2
0
9 2-In AND~
219 698 635 0 3 22
0 20 23 14
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U3D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
659 0 0
2
43239.8 1
0
9 2-In AND~
219 698 598 0 3 22
0 20 21 13
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U3C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3800 0 0
2
43239.8 0
0
7 Ground~
168 413 735 0 1 3
0 2
0
0 0 53360 270
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6792 0 0
2
43239.8 0
0
7 Ground~
168 408 647 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3701 0 0
2
43239.8 0
0
2 +V
167 393 684 0 1 3
0 24
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V6
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6316 0 0
2
43239.8 0
0
7 74LS283
152 451 691 0 14 29
0 2 2 2 24 25 26 27 28 2
21 23 19 22 51
0
0 0 4336 0
7 74LS283
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
8734 0 0
2
43239.8 0
0
7 Ground~
168 597 198 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7988 0 0
2
43239.7 0
0
9 2-In AND~
219 353 626 0 3 22
0 25 26 30
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U3B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3217 0 0
2
43239.7 0
0
7 74LS293
154 296 673 0 8 17
0 30 30 17 28 25 26 27 28
0
0 0 4336 0
7 74LS293
-24 -35 25 -27
2 U6
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 0 0 0 0
1 U
3965 0 0
2
43239.7 0
0
7 74LS151
20 542 244 0 14 29
0 52 53 54 55 43 44 45 46 2
2 32 31 56 8
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
8239 0 0
2
43239.7 0
0
7 74LS293
154 339 526 0 8 17
0 29 29 33 31 57 29 32 31
0
0 0 4336 0
7 74LS293
-24 -35 25 -27
2 U4
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 0 0 0 0
1 U
828 0 0
2
43239.7 0
0
9 2-In AND~
219 204 598 0 3 22
0 33 37 38
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6187 0 0
2
43239.7 0
0
7 74LS293
154 170 526 0 8 17
0 38 38 17 37 58 59 33 37
0
0 0 4336 0
7 74LS293
-24 -35 25 -27
2 U2
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 0 0 0 0
1 U
7107 0 0
2
43239.7 0
0
7 Pulser~
4 101 827 0 10 12
0 60 61 18 62 0 0 10 10 6
7
0
0 0 4144 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6433 0 0
2
43239.7 0
0
7 Ground~
168 93 409 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8559 0 0
2
43239.7 0
0
7 74LS139
118 142 393 0 14 29
0 33 37 2 63 64 65 66 34 35
36 67 68 69 70
0
0 0 4336 0
7 74LS139
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 0 0 0 0
1 U
3674 0 0
2
43239.7 0
0
2 +V
167 117 299 0 1 3
0 39
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V4
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5697 0 0
2
43239.7 0
0
2 +V
167 118 233 0 1 3
0 40
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3805 0 0
2
43239.7 0
0
2 +V
167 118 171 0 1 3
0 41
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5219 0 0
2
43239.7 0
0
2 +V
167 118 113 0 1 3
0 42
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3795 0 0
2
43239.7 0
0
14 NO PushButton~
191 217 274 0 2 5
0 43 36
0
0 0 4720 0
0
3 AST
-9 -21 12 -13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3637 0 0
2
43239.7 2
0
14 NO PushButton~
191 316 274 0 2 5
0 43 35
0
0 0 4720 0
0
2 b0
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3226 0 0
2
43239.7 1
0
14 NO PushButton~
191 419 274 0 2 5
0 43 34
0
0 0 4720 0
0
6 TRALHA
-15 -20 27 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
6966 0 0
2
43239.7 0
0
14 NO PushButton~
191 217 208 0 2 5
0 44 36
0
0 0 4720 0
0
2 b7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
9796 0 0
2
43239.7 2
0
14 NO PushButton~
191 316 208 0 2 5
0 44 35
0
0 0 4720 0
0
2 b8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
5952 0 0
2
43239.7 1
0
14 NO PushButton~
191 419 208 0 2 5
0 44 34
0
0 0 4720 0
0
2 b9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3649 0 0
2
43239.7 0
0
14 NO PushButton~
191 217 146 0 2 5
0 45 36
0
0 0 4720 0
0
2 b4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3716 0 0
2
43239.7 2
0
14 NO PushButton~
191 316 146 0 2 5
0 45 35
0
0 0 4720 0
0
2 b5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4797 0 0
2
43239.7 1
0
14 NO PushButton~
191 419 146 0 2 5
0 45 34
0
0 0 4720 0
0
2 b6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4681 0 0
2
43239.7 0
0
14 NO PushButton~
191 418 88 0 2 5
0 46 34
0
0 0 4720 0
0
2 b3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
9730 0 0
2
43239.7 0
0
14 NO PushButton~
191 315 88 0 2 5
0 46 35
0
0 0 4720 0
0
2 b2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
9874 0 0
2
43239.7 0
0
14 NO PushButton~
191 216 88 0 2 5
0 46 36
0
0 0 4720 0
0
2 b1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
364 0 0
2
43239.7 0
0
9 Resistor~
219 145 297 0 3 5
0 39 43 1
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 266
82 0 0 0 1 0 0 0
1 R
3656 0 0
2
43239.7 0
0
9 Resistor~
219 146 231 0 3 5
0 40 44 1
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 250
82 0 0 0 1 0 0 0
1 R
3131 0 0
2
43239.7 0
0
9 Resistor~
219 146 169 0 3 5
0 41 45 1
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 38
82 0 0 0 1 0 0 0
1 R
6772 0 0
2
43239.7 0
0
9 Resistor~
219 146 111 0 3 5
0 42 46 1
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 26
82 0 0 0 1 0 0 0
1 R
9557 0 0
2
43239.7 0
0
91
2 2 3 0 0 4224 0 2 7 0 0 4
710 562
748 562
748 550
785 550
2 1 4 0 0 4224 0 3 2 0 0 2
666 562
674 562
2 1 5 0 0 4224 0 4 3 0 0 2
623 562
630 562
2 1 6 0 0 4224 0 5 4 0 0 2
576 562
587 562
1 1 7 0 0 8320 0 7 1 0 0 3
779 541
773 541
773 455
0 1 8 0 0 4096 0 0 5 40 0 2
510 562
540 562
7 4 9 0 0 4224 0 7 6 0 0 3
849 541
888 541
888 509
9 3 10 0 0 8320 0 7 6 0 0 3
849 559
894 559
894 509
11 2 11 0 0 8320 0 7 6 0 0 3
849 577
900 577
900 509
13 1 12 0 0 8320 0 7 6 0 0 3
849 595
906 595
906 509
3 3 13 0 0 4224 0 13 7 0 0 4
719 598
758 598
758 568
785 568
3 4 14 0 0 8320 0 12 7 0 0 4
719 635
765 635
765 577
785 577
3 5 15 0 0 8320 0 10 7 0 0 4
719 672
772 672
772 586
785 586
3 6 16 0 0 8320 0 9 7 0 0 4
719 708
780 708
780 595
785 595
3 0 17 0 0 4096 0 8 0 0 70 2
165 720
165 682
3 1 18 0 0 8320 0 25 8 0 0 3
125 818
156 818
156 766
2 0 19 0 0 4096 0 11 0 0 26 2
591 668
591 700
1 0 20 0 0 4096 0 12 0 0 20 2
674 626
661 626
1 0 20 0 0 0 0 10 0 0 20 2
674 663
661 663
0 1 20 0 0 4224 0 0 9 21 0 3
661 589
661 699
674 699
4 1 20 0 0 0 0 11 13 0 0 3
591 617
591 589
674 589
3 0 21 0 0 4096 0 11 0 0 24 2
600 668
600 682
1 0 22 0 0 4096 0 11 0 0 27 2
582 668
582 709
10 2 21 0 0 4224 0 17 13 0 0 4
483 682
630 682
630 607
674 607
11 2 23 0 0 4224 0 17 12 0 0 4
483 691
639 691
639 644
674 644
12 2 19 0 0 4224 0 17 10 0 0 4
483 700
647 700
647 681
674 681
13 2 22 0 0 4224 0 17 9 0 0 4
483 709
631 709
631 717
674 717
1 9 2 0 0 4096 0 14 17 0 0 2
420 736
419 736
1 0 2 0 0 0 0 15 0 0 30 2
408 655
408 655
1 0 2 0 0 4096 0 17 0 0 31 3
419 655
408 655
408 664
3 2 2 0 0 0 0 17 17 0 0 4
419 673
408 673
408 664
419 664
1 4 24 0 0 4224 0 16 17 0 0 2
404 682
419 682
0 5 25 0 0 12416 0 0 17 44 0 4
342 664
348 664
348 691
419 691
0 6 26 0 0 8320 0 0 17 43 0 3
342 673
342 700
419 700
7 7 27 0 0 12416 0 20 17 0 0 4
328 682
338 682
338 709
419 709
8 8 28 0 0 12416 0 20 17 0 0 4
328 691
334 691
334 718
419 718
10 0 2 0 0 4224 0 21 0 0 39 3
574 226
597 226
597 217
6 0 29 0 0 12416 0 22 0 0 48 5
371 526
381 526
381 565
295 565
295 526
9 1 2 0 0 128 0 21 18 0 0 3
580 217
597 217
597 206
14 2 8 0 0 12416 0 21 8 0 0 6
580 280
580 304
510 304
510 788
174 788
174 766
2 0 30 0 0 4096 0 20 0 0 42 3
264 673
252 673
252 664
3 1 30 0 0 4224 0 19 20 0 0 4
352 602
252 602
252 664
264 664
6 2 26 0 0 0 0 20 19 0 0 3
328 673
361 673
361 647
5 1 25 0 0 0 0 20 19 0 0 3
328 664
343 664
343 647
4 8 28 0 0 0 0 20 20 0 0 4
258 691
258 708
328 708
328 691
8 12 31 0 0 8320 0 22 21 0 0 4
371 544
596 544
596 244
574 244
7 11 32 0 0 8320 0 22 21 0 0 4
371 535
606 535
606 235
574 235
2 1 29 0 0 0 0 22 22 0 0 4
307 526
295 526
295 517
307 517
4 8 31 0 0 0 0 22 22 0 0 4
301 544
301 558
371 558
371 544
0 3 33 0 0 8192 0 0 22 63 0 3
211 536
211 535
301 535
2 2 34 0 0 8192 0 40 41 0 0 3
402 154
401 154
401 96
2 2 34 0 0 4096 0 37 40 0 0 2
402 216
402 154
2 2 34 0 0 4096 0 34 37 0 0 2
402 282
402 216
8 2 34 0 0 4224 0 27 34 0 0 3
180 375
402 375
402 282
2 2 35 0 0 8192 0 39 42 0 0 3
299 154
298 154
298 96
2 2 35 0 0 4096 0 36 39 0 0 2
299 216
299 154
2 2 35 0 0 4096 0 33 36 0 0 2
299 282
299 216
9 2 35 0 0 4224 0 27 33 0 0 3
180 384
299 384
299 282
2 2 36 0 0 8192 0 38 43 0 0 3
200 154
199 154
199 96
2 2 36 0 0 4096 0 35 38 0 0 2
200 216
200 154
2 2 36 0 0 4096 0 32 35 0 0 2
200 282
200 216
10 2 36 0 0 8320 0 27 32 0 0 3
180 393
200 393
200 282
0 1 33 0 0 8320 0 0 27 68 0 5
211 537
211 465
68 465
68 375
110 375
8 2 37 0 0 12416 0 24 27 0 0 6
202 544
226 544
226 455
76 455
76 384
110 384
2 0 38 0 0 4096 0 24 0 0 66 2
138 526
126 526
3 1 38 0 0 8320 0 23 24 0 0 4
202 621
126 621
126 517
138 517
2 0 37 0 0 0 0 23 0 0 69 2
193 576
193 560
1 7 33 0 0 0 0 23 24 0 0 3
211 576
211 535
202 535
8 4 37 0 0 0 0 24 24 0 0 4
202 544
202 560
132 560
132 544
3 3 17 0 0 4224 0 20 24 0 0 4
258 682
87 682
87 535
132 535
1 3 2 0 0 128 0 26 27 0 0 3
93 403
93 393
104 393
1 1 39 0 0 4224 0 28 44 0 0 2
128 297
127 297
1 1 40 0 0 4224 0 29 45 0 0 2
129 231
128 231
1 1 41 0 0 4224 0 30 46 0 0 2
129 169
128 169
1 1 42 0 0 4224 0 31 47 0 0 2
129 111
128 111
1 0 43 0 0 4096 0 34 0 0 79 2
436 282
436 297
1 0 43 0 0 0 0 33 0 0 79 2
333 282
333 297
1 0 43 0 0 0 0 32 0 0 79 2
234 282
234 297
2 5 43 0 0 4224 0 44 21 0 0 4
163 297
481 297
481 253
510 253
1 0 44 0 0 4096 0 37 0 0 83 2
436 216
436 231
1 0 44 0 0 0 0 36 0 0 83 2
333 216
333 231
1 0 44 0 0 0 0 35 0 0 83 2
234 216
234 231
2 6 44 0 0 4224 0 45 21 0 0 4
164 231
488 231
488 262
510 262
1 0 45 0 0 4096 0 40 0 0 87 2
436 154
436 169
1 0 45 0 0 0 0 39 0 0 87 2
333 154
333 169
1 0 45 0 0 0 0 38 0 0 87 2
234 154
234 169
2 7 45 0 0 4224 0 46 21 0 0 4
164 169
496 169
496 271
510 271
1 0 46 0 0 4096 0 41 0 0 91 2
435 96
435 111
1 0 46 0 0 0 0 42 0 0 91 2
332 96
332 111
1 0 46 0 0 0 0 43 0 0 91 2
233 96
233 111
2 8 46 0 0 4224 0 47 21 0 0 4
164 111
503 111
503 280
510 280
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
