CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 26 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
35
7 74LS165
97 455 231 0 14 29
0 59 60 61 62 55 56 57 58 29
6 2 7 73 28
0
0 0 4320 0
7 74LS165
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 1 0 0
1 U
5130 0 0
2
43198.6 34
0
8 Hex Key~
166 410 177 0 11 12
0 58 57 56 55 0 0 0 0 0
2 50
0
0 0 4128 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
391 0 0
2
43198.6 33
0
8 Hex Key~
166 372 177 0 11 12
0 62 61 60 59 0 0 0 0 0
4 52
0
0 0 4128 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3124 0 0
2
43198.6 32
0
7 Ground~
168 508 245 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
43198.6 31
0
7 Ground~
168 335 250 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
43198.6 30
0
8 Hex Key~
166 199 182 0 11 12
0 54 53 52 51 0 0 0 0 0
2 50
0
0 0 4128 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5572 0 0
2
43198.6 29
0
8 Hex Key~
166 237 182 0 11 12
0 50 49 48 47 0 0 0 0 0
4 52
0
0 0 4128 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8901 0 0
2
43198.6 28
0
7 74LS165
97 282 236 0 14 29
0 51 52 53 54 47 48 49 50 30
6 2 7 72 29
0
0 0 4320 0
7 74LS165
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 1 0 0
1 U
7361 0 0
2
43198.6 27
0
7 Ground~
168 159 253 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
43198.6 26
0
8 Hex Key~
166 23 185 0 11 12
0 46 45 44 43 0 0 0 0 0
1 49
0
0 0 4128 0
0
4 KPD5
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
972 0 0
2
43198.6 25
0
8 Hex Key~
166 61 185 0 11 12
0 42 41 40 39 0 0 0 0 0
8 56
0
0 0 4128 0
0
4 KPD6
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3472 0 0
2
43198.6 24
0
7 74LS165
97 106 239 0 14 29
0 43 44 45 46 39 40 41 42 26
6 2 7 71 30
0
0 0 4320 0
7 74LS165
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 1 0 0
1 U
9998 0 0
2
43198.6 23
0
7 Ground~
168 696 244 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
43198.6 22
0
8 Hex Key~
166 560 176 0 11 12
0 38 37 36 35 0 0 0 0 0
8 56
0
0 0 4128 0
0
4 KPD7
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4597 0 0
2
43198.6 21
0
8 Hex Key~
166 598 176 0 11 12
0 34 33 32 31 0 0 0 0 0
1 49
0
0 0 4128 0
0
4 KPD8
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3835 0 0
2
43198.6 20
0
7 74LS165
97 643 230 0 14 29
0 35 36 37 38 31 32 33 34 28
6 2 7 70 26
0
0 0 4320 0
7 74LS165
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 1 0 0
1 U
3670 0 0
2
43198.6 19
0
7 74LS164
127 756 252 0 12 25
0 26 26 7 27 25 23 22 21 20
19 18 17
0
0 0 4320 0
7 74LS164
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
5616 0 0
2
43198.6 18
0
2 +V
167 710 296 0 1 3
0 27
0
0 0 61664 180
2 5V
7 -2 21 6
2 V2
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
43198.6 17
0
7 74LS293
154 726 64 0 8 17
0 2 2 2 7 3 67 68 69
0
0 0 4832 512
7 74LS293
-24 -35 25 -27
4 Div8
-20 -36 8 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
43198.6 16
0
7 Ground~
168 777 55 0 1 3
0 2
0
0 0 53344 90
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
43198.6 15
0
7 74LS273
150 854 243 0 18 37
0 24 5 25 23 22 21 20 19 18
17 16 15 14 13 9 10 11 12
0
0 0 4320 0
7 74LS273
-24 -60 25 -52
2 U7
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
4299 0 0
2
43198.6 14
0
2 +V
167 811 187 0 1 3
0 24
0
0 0 61664 512
2 5V
7 -2 21 6
2 V1
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
43198.6 13
0
14 Logic Display~
6 938 188 0 1 2
10 16
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R8
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
43198.6 12
0
14 Logic Display~
6 938 208 0 1 2
10 15
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R7
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
43198.6 11
0
14 Logic Display~
6 938 229 0 1 2
10 14
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R6
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
43198.6 10
0
14 Logic Display~
6 939 250 0 1 2
10 13
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R5
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
43198.6 9
0
14 Logic Display~
6 940 270 0 1 2
10 9
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R4
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
43198.6 8
0
14 Logic Display~
6 940 291 0 1 2
10 10
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R3
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
43198.6 7
0
14 Logic Display~
6 940 314 0 1 2
10 11
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R2
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
43198.6 6
0
14 Logic Display~
6 940 338 0 1 2
10 12
0
0 0 53344 270
6 100MEG
3 -16 45 -8
2 R1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
43198.6 5
0
7 Pulser~
4 822 138 0 10 12
0 64 65 7 66 0 0 10 10 2
8
0
0 0 4640 512
0
5 Clock
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3409 0 0
2
43198.6 4
0
5 7474~
219 578 91 0 6 22
0 8 3 7 8 63 4
0
0 0 4192 512
4 7474
7 -60 35 -52
3 U5A
27 -61 48 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3951 0 0
2
43198.6 3
0
2 +V
167 618 19 0 1 3
0 8
0
0 0 61664 512
2 5V
7 -2 21 6
2 V4
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8885 0 0
2
43198.6 2
0
8 2-In OR~
219 371 91 0 3 22
0 6 7 6
0
0 0 96 90
6 74LS32
-21 -24 21 -16
3 U9A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3780 0 0
2
43198.6 1
0
9 Inverter~
13 658 113 0 2 22
0 4 5
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
9265 0 0
2
43198.6 0
0
82
2 5 3 0 0 16 0 32 19 0 0 2
608 55
688 55
1 6 4 0 0 16 0 35 32 0 0 4
643 113
551 113
551 55
560 55
2 2 5 0 0 16 0 35 21 0 0 6
679 113
745 113
745 168
790 168
790 216
822 216
3 0 6 0 0 16 0 34 0 0 42 3
374 61
400 61
400 125
2 0 7 0 0 16 0 34 0 0 40 2
383 107
383 140
1 3 6 0 0 16 0 34 34 0 0 5
365 107
365 117
349 117
349 61
374 61
1 0 8 0 0 16 0 33 0 0 8 2
618 28
618 28
4 1 8 0 0 16 0 32 32 0 0 4
584 103
618 103
618 28
584 28
3 0 7 0 0 16 0 32 0 0 28 2
608 73
608 140
15 1 9 0 0 16 0 21 27 0 0 4
886 261
909 261
909 274
924 274
16 1 10 0 0 16 0 21 28 0 0 4
886 270
899 270
899 295
924 295
17 1 11 0 0 16 0 21 29 0 0 4
886 279
892 279
892 318
924 318
18 1 12 0 0 16 0 21 30 0 0 3
886 288
886 342
924 342
14 1 13 0 0 16 0 21 26 0 0 3
886 252
886 254
923 254
13 1 14 0 0 16 0 21 25 0 0 4
886 243
895 243
895 233
922 233
1 12 15 0 0 16 0 24 21 0 0 4
922 212
891 212
891 234
886 234
11 1 16 0 0 16 0 21 23 0 0 3
886 225
886 192
922 192
12 10 17 0 0 16 0 17 21 0 0 2
788 288
822 288
11 9 18 0 0 16 0 17 21 0 0 2
788 279
822 279
10 8 19 0 0 16 0 17 21 0 0 2
788 270
822 270
9 7 20 0 0 16 0 17 21 0 0 2
788 261
822 261
8 6 21 0 0 16 0 17 21 0 0 2
788 252
822 252
7 5 22 0 0 16 0 17 21 0 0 2
788 243
822 243
6 4 23 0 0 16 0 17 21 0 0 2
788 234
822 234
1 1 24 0 0 16 0 21 22 0 0 3
816 207
811 207
811 196
5 3 25 0 0 16 0 17 21 0 0 2
788 225
822 225
0 0 7 0 0 16 0 0 0 32 33 2
688 140
716 140
0 12 7 0 0 16 0 0 1 0 0 4
652 140
502 140
502 222
487 222
0 1 2 0 0 16 0 0 20 30 0 2
758 56
770 56
3 1 2 0 0 16 0 19 19 0 0 3
758 73
758 55
752 55
2 1 2 0 0 16 0 19 19 0 0 2
752 64
752 55
12 0 7 0 0 16 0 16 0 0 28 4
675 221
688 221
688 140
652 140
3 3 7 0 0 16 0 31 17 0 0 4
798 129
716 129
716 252
724 252
0 4 7 0 0 16 0 0 19 33 0 3
781 129
781 82
758 82
0 1 26 0 0 16 0 0 17 38 0 4
679 266
707 266
707 225
724 225
1 4 27 0 0 16 0 18 17 0 0 3
710 281
710 270
718 270
2 1 26 0 0 16 0 17 17 0 0 2
724 234
724 225
14 9 26 0 0 16 0 16 12 0 0 6
675 266
679 266
679 293
147 293
147 203
138 203
12 0 7 0 0 16 0 12 0 0 40 4
138 230
152 230
152 140
328 140
12 0 7 0 0 16 0 8 0 0 28 4
314 227
328 227
328 140
502 140
10 0 6 0 0 16 0 12 0 0 42 3
144 212
144 125
320 125
10 0 6 0 0 16 0 8 0 0 43 3
320 209
320 125
493 125
10 10 6 0 0 16 0 1 16 0 0 4
493 204
493 125
681 125
681 203
14 9 28 0 0 16 0 1 16 0 0 5
487 267
538 267
538 146
675 146
675 194
14 9 29 0 0 16 0 8 1 0 0 5
314 272
350 272
350 148
487 148
487 195
14 9 30 0 0 16 0 12 8 0 0 5
138 275
175 275
175 153
314 153
314 200
1 11 2 0 0 16 0 13 16 0 0 3
696 238
696 212
681 212
5 4 31 0 0 16 0 16 15 0 0 3
611 239
589 239
589 200
6 3 32 0 0 16 0 16 15 0 0 3
611 248
595 248
595 200
2 7 33 0 0 16 0 15 16 0 0 3
601 200
601 257
611 257
1 8 34 0 0 16 0 15 16 0 0 3
607 200
607 266
611 266
1 4 35 0 0 16 0 16 14 0 0 3
611 203
551 203
551 200
3 2 36 0 0 16 0 14 16 0 0 3
557 200
557 212
611 212
3 2 37 0 0 16 0 16 14 0 0 3
611 221
563 221
563 200
1 4 38 0 0 16 0 14 16 0 0 3
569 200
569 230
611 230
1 11 2 0 0 16 0 9 12 0 0 3
159 247
159 221
144 221
5 4 39 0 0 16 0 12 11 0 0 3
74 248
52 248
52 209
6 3 40 0 0 16 0 12 11 0 0 3
74 257
58 257
58 209
2 7 41 0 0 16 0 11 12 0 0 3
64 209
64 266
74 266
1 8 42 0 0 16 0 11 12 0 0 3
70 209
70 275
74 275
1 4 43 0 0 16 0 12 10 0 0 3
74 212
14 212
14 209
3 2 44 0 0 16 0 10 12 0 0 3
20 209
20 221
74 221
3 2 45 0 0 16 0 12 10 0 0 3
74 230
26 230
26 209
1 4 46 0 0 16 0 10 12 0 0 3
32 209
32 239
74 239
1 11 2 0 0 16 0 5 8 0 0 3
335 244
335 218
320 218
5 4 47 0 0 16 0 8 7 0 0 3
250 245
228 245
228 206
6 3 48 0 0 16 0 8 7 0 0 3
250 254
234 254
234 206
2 7 49 0 0 16 0 7 8 0 0 3
240 206
240 263
250 263
1 8 50 0 0 16 0 7 8 0 0 3
246 206
246 272
250 272
1 4 51 0 0 16 0 8 6 0 0 3
250 209
190 209
190 206
3 2 52 0 0 16 0 6 8 0 0 3
196 206
196 218
250 218
3 2 53 0 0 16 0 8 6 0 0 3
250 227
202 227
202 206
1 4 54 0 0 16 0 6 8 0 0 3
208 206
208 236
250 236
1 11 2 0 0 16 0 4 1 0 0 3
508 239
508 213
493 213
5 4 55 0 0 16 0 1 2 0 0 3
423 240
401 240
401 201
6 3 56 0 0 16 0 1 2 0 0 3
423 249
407 249
407 201
2 7 57 0 0 16 0 2 1 0 0 3
413 201
413 258
423 258
1 8 58 0 0 16 0 2 1 0 0 3
419 201
419 267
423 267
1 4 59 0 0 16 0 1 3 0 0 3
423 204
363 204
363 201
3 2 60 0 0 16 0 3 1 0 0 3
369 201
369 213
423 213
3 2 61 0 0 16 0 1 3 0 0 3
423 222
375 222
375 201
1 4 62 0 0 16 0 3 1 0 0 3
381 201
381 231
423 231
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
