CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 170 30 100 10
1131 88 1917 1018
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
1299 184 1412 281
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 259 917 0 1 11
0 15
0
0 0 21360 90
2 0V
11 0 25 8
1 D
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
361 0 0
2
43185 0
0
13 Logic Switch~
5 194 917 0 1 11
0 22
0
0 0 21360 90
2 0V
11 0 25 8
1 C
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3343 0 0
2
43185 0
0
13 Logic Switch~
5 129 919 0 1 11
0 16
0
0 0 21360 90
2 0V
11 0 25 8
1 B
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7923 0 0
2
43185 0
0
13 Logic Switch~
5 71 919 0 1 11
0 21
0
0 0 21360 90
2 0V
11 0 25 8
1 A
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6174 0 0
2
43185 0
0
14 Logic Display~
6 547 705 0 1 2
10 2
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S0
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6692 0 0
2
43185 0
0
14 Logic Display~
6 552 566 0 1 2
10 3
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8790 0 0
2
43185 0
0
14 Logic Display~
6 550 442 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4595 0 0
2
43185 0
0
14 Logic Display~
6 556 330 0 1 2
10 5
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 S3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
667 0 0
2
43185 0
0
5 4071~
219 483 710 0 3 22
0 7 6 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
8743 0 0
2
43185 0
0
5 4071~
219 477 447 0 3 22
0 12 11 4
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
8298 0 0
2
43185 0
0
5 4071~
219 489 335 0 3 22
0 14 13 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
313 0 0
2
43185 0
0
8 3-In OR~
219 486 571 0 4 22
0 10 9 8 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
7548 0 0
2
43185 0
0
9 Inverter~
13 277 844 0 2 22
0 15 18
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
8973 0 0
2
43185 0
0
9 Inverter~
13 212 843 0 2 22
0 22 20
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
9712 0 0
2
43185 0
0
9 Inverter~
13 150 845 0 2 22
0 16 19
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
4518 0 0
2
43185 0
0
9 Inverter~
13 88 846 0 2 22
0 21 17
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
5596 0 0
2
43185 0
0
9 2-In AND~
219 416 684 0 3 22
0 19 18 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
692 0 0
2
43185 1
0
9 3-In AND~
219 414 741 0 4 22
0 17 16 15 6
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 3 0
1 U
6258 0 0
2
43185 0
0
9 3-In AND~
219 417 526 0 4 22
0 17 19 15 10
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
5578 0 0
2
43185 0
0
9 3-In AND~
219 414 634 0 4 22
0 21 20 18 8
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 1 0
1 U
8709 0 0
2
43185 1
0
9 2-In AND~
219 416 577 0 3 22
0 17 22 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9131 0 0
2
43185 0
0
9 3-In AND~
219 416 481 0 4 22
0 21 20 18 11
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
3645 0 0
2
43185 1
0
9 2-In AND~
219 414 421 0 3 22
0 17 16 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7613 0 0
2
43185 0
0
9 2-In AND~
219 414 306 0 3 22
0 21 22 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9467 0 0
2
43185 0
0
9 3-In AND~
219 416 366 0 4 22
0 21 19 15 13
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
3932 0 0
2
43185 0
0
48
3 1 2 0 0 4224 0 9 5 0 0 4
516 710
524 710
524 709
531 709
4 1 3 0 0 4224 0 12 6 0 0 4
519 571
529 571
529 570
536 570
3 1 4 0 0 4224 0 10 7 0 0 4
510 447
527 447
527 446
534 446
3 1 5 0 0 4224 0 11 8 0 0 4
522 335
533 335
533 334
540 334
4 2 6 0 0 4224 0 18 9 0 0 4
435 741
462 741
462 719
470 719
3 1 7 0 0 4224 0 17 9 0 0 4
437 684
462 684
462 701
470 701
4 3 8 0 0 8320 0 20 12 0 0 4
435 634
465 634
465 580
473 580
3 2 9 0 0 4224 0 21 12 0 0 4
437 577
465 577
465 571
474 571
4 1 10 0 0 8320 0 19 12 0 0 4
438 526
465 526
465 562
473 562
4 2 11 0 0 8320 0 22 10 0 0 4
437 481
456 481
456 456
464 456
3 1 12 0 0 4224 0 23 10 0 0 4
435 421
456 421
456 438
464 438
4 2 13 0 0 4224 0 25 11 0 0 4
437 366
468 366
468 344
476 344
3 1 14 0 0 4224 0 24 11 0 0 4
435 306
468 306
468 326
476 326
3 0 15 0 0 4096 0 18 0 0 38 2
390 750
260 750
2 0 16 0 0 4096 0 18 0 0 42 2
390 741
130 741
1 0 17 0 0 4096 0 18 0 0 44 2
390 732
91 732
2 0 18 0 0 4096 0 17 0 0 39 2
392 693
280 693
1 0 19 0 0 4096 0 17 0 0 43 2
392 675
153 675
3 0 18 0 0 0 0 20 0 0 39 2
390 643
280 643
2 0 20 0 0 4096 0 20 0 0 40 2
390 634
215 634
1 0 21 0 0 4096 0 20 0 0 37 2
390 625
72 625
2 0 22 0 0 4096 0 21 0 0 41 2
392 586
195 586
1 0 17 0 0 4096 0 21 0 0 44 2
392 568
91 568
3 0 15 0 0 4096 0 19 0 0 38 2
393 535
260 535
2 0 19 0 0 4096 0 19 0 0 43 2
393 526
153 526
1 0 17 0 0 4096 0 19 0 0 44 2
393 517
91 517
3 0 18 0 0 0 0 22 0 0 39 2
392 490
280 490
2 0 20 0 0 4096 0 22 0 0 40 2
392 481
215 481
1 0 21 0 0 4096 0 22 0 0 37 2
392 472
72 472
2 0 16 0 0 0 0 23 0 0 42 2
390 430
130 430
1 0 17 0 0 0 0 23 0 0 44 2
390 412
91 412
3 0 15 0 0 0 0 25 0 0 38 2
392 375
260 375
2 0 19 0 0 0 0 25 0 0 43 2
392 366
153 366
1 0 21 0 0 0 0 25 0 0 37 2
392 357
72 357
2 0 22 0 0 0 0 24 0 0 41 2
390 315
195 315
1 0 21 0 0 0 0 24 0 0 37 2
390 297
72 297
0 0 21 0 0 4224 0 0 0 48 0 2
72 866
72 216
0 0 15 0 0 4224 0 0 0 45 0 2
260 862
260 218
2 0 18 0 0 4224 0 13 0 0 0 2
280 826
280 219
2 0 20 0 0 4224 0 14 0 0 0 2
215 825
215 218
0 0 22 0 0 4224 0 0 0 46 0 2
195 861
195 217
0 0 16 0 0 4224 0 0 0 47 0 2
130 864
130 216
2 0 19 0 0 4224 0 15 0 0 0 2
153 827
153 217
2 0 17 0 0 4224 0 16 0 0 0 2
91 828
91 216
1 1 15 0 0 0 0 1 13 0 0 3
260 904
260 862
280 862
1 1 22 0 0 0 0 2 14 0 0 3
195 904
195 861
215 861
1 1 16 0 0 0 0 3 15 0 0 3
130 906
130 863
153 863
1 1 21 0 0 0 0 4 16 0 0 3
72 906
72 864
91 864
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
