CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
39
8 2-In OR~
219 782 437 0 3 22
0 3 4 4
0
0 0 112 90
6 74LS32
-21 -24 21 -16
3 U7A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8464 0 0
2
5.89842e-315 0
0
7 Output~
178 829 508 0 17 19
0 3 0 0 0 0 0 0 0 0
67 108 111 99 107 32 32 32
0
0 0 53360 0
0
2 T2
-13 -26 1 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7168 0 0
2
5.89842e-315 0
0
6 Input~
177 271 85 0 17 19
0 3 0 0 0 0 0 0 0 0
67 108 111 99 107 32 32 32
0
0 0 53360 0
0
2 T1
-7 -26 7 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3171 0 0
2
5.89842e-315 0
0
9 Inverter~
13 672 272 0 2 22
0 7 6
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4139 0 0
2
5.89842e-315 0
0
5 7474~
219 785 345 0 6 22
0 6 2 2 4 53 5
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U4A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
6435 0 0
2
5.89842e-315 5.30499e-315
0
7 Ground~
168 753 333 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5283 0 0
2
5.89842e-315 5.26354e-315
0
2 +V
167 495 136 0 1 3
0 12
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V6
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6874 0 0
2
5.89842e-315 0
0
7 Ground~
168 505 187 0 1 3
0 2
0
0 0 53360 270
0
5 GND12
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5305 0 0
2
5.89842e-315 0
0
7 74LS283
152 551 143 0 14 29
0 2 2 2 12 2 2 13 14 2
8 9 10 11 54
0
0 0 4336 0
7 74LS283
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.89842e-315 0
0
14 Logic Display~
6 854 182 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
6 ALARME
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
43205.8 0
0
7 Ground~
168 680 196 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8402 0 0
2
43205.8 1
0
12 Hex Display~
7 726 155 0 16 19
10 18 17 16 15 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
4 Temp
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3751 0 0
2
43205.8 2
0
12 Hex Display~
7 689 155 0 16 19
10 19 2 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 Temp
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4292 0 0
2
43205.8 3
0
7 Ground~
168 606 416 0 1 3
0 2
0
0 0 53360 270
0
5 GND10
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6118 0 0
2
43205.8 4
0
7 74LS283
152 665 372 0 14 29
0 24 23 22 21 2 20 20 2 2
15 16 17 18 19
0
0 0 4336 0
7 74LS283
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
43205.8 5
0
7 Ground~
168 642 494 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
43205.8 6
0
7 Ground~
168 641 251 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
319 0 0
2
43205.8 7
0
7 Ground~
168 552 523 0 1 3
0 2
0
0 0 53360 270
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3976 0 0
2
43205.8 8
0
2 +V
167 557 508 0 1 3
0 25
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V4
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7634 0 0
2
43205.8 9
0
6 74LS85
106 606 497 0 14 29
0 24 23 22 21 25 2 2 25 2
26 2 55 56 20
0
0 0 4336 0
6 74LS85
-21 -52 21 -44
2 U2
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
523 0 0
2
43205.8 10
0
2 +V
167 659 480 0 1 3
0 26
0
0 0 53616 270
2 5V
-7 -15 7 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6748 0 0
2
43205.8 11
0
2 +V
167 658 237 0 1 3
0 27
0
0 0 53616 270
2 5V
-7 -15 7 -7
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6901 0 0
2
43205.8 12
0
2 +V
167 546 229 0 1 3
0 28
0
0 0 53616 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
842 0 0
2
43205.8 13
0
7 Ground~
168 534 235 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3277 0 0
2
43205.8 14
0
6 74LS85
106 603 254 0 14 29
0 28 2 28 28 24 23 22 21 2
27 2 7 57 58
0
0 0 4336 0
6 74LS85
-21 -52 21 -44
2 U1
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4212 0 0
2
43205.8 15
0
12 Hex Display~
7 635 113 0 16 19
10 11 10 9 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
6 Tanque
-21 -38 21 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4720 0 0
2
43205.8 16
0
7 Pulser~
4 255 140 0 10 12
0 59 60 3 61 0 0 10 10 11
7
0
0 0 4656 0
0
5 Clock
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5551 0 0
2
43205.8 17
0
7 Ground~
168 337 179 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6986 0 0
2
43205.8 18
0
7 74LS293
154 383 139 0 8 17
0 2 2 2 3 62 13 14 63
0
0 0 4848 0
0
4 Div4
-14 -36 14 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
8745 0 0
2
43205.8 19
0
7 Ground~
168 361 557 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9592 0 0
2
43205.8 20
0
7 Ground~
168 361 353 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8748 0 0
2
43205.8 21
0
7 Ground~
168 487 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
43205.8 22
0
7 74LS157
122 515 383 0 14 29
0 13 48 49 47 50 46 51 45 52
2 24 23 22 21
0
0 0 4336 0
7 74LS157
-24 -60 25 -52
2 A1
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
631 0 0
2
43205.8 23
0
7 74LS157
122 399 491 0 14 29
0 14 29 33 30 34 31 35 32 36
2 48 47 46 45
0
0 0 4336 0
7 74LS157
-24 -60 25 -52
2 A2
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9466 0 0
2
43205.8 24
0
7 74LS157
122 399 288 0 14 29
0 14 37 41 38 42 39 43 40 44
2 49 50 51 52
0
0 0 4336 0
7 74LS157
-24 -60 25 -52
2 A3
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3266 0 0
2
43205.8 25
0
8 Hex Key~
166 219 524 0 11 12
0 32 31 30 29 0 0 0 0 0
12 67
0
0 0 4656 0
0
7 Tanque3
-24 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7693 0 0
2
43205.8 26
0
8 Hex Key~
166 218 420 0 11 12
0 36 35 34 33 0 0 0 0 0
0 48
0
0 0 4656 0
0
7 Tanque2
-24 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3723 0 0
2
43205.8 27
0
8 Hex Key~
166 219 322 0 11 12
0 40 39 38 37 0 0 0 0 0
9 57
0
0 0 4656 0
0
7 Tanque1
-24 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3440 0 0
2
43205.8 28
0
8 Hex Key~
166 220 222 0 11 12
0 44 43 42 41 0 0 0 0 0
11 66
0
0 0 4656 0
0
7 Tanque0
-24 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6263 0 0
2
43205.8 29
0
95
2 0 4 0 0 12416 0 1 0 0 2 5
794 453
794 464
809 464
809 395
785 395
3 4 4 0 0 0 0 1 5 0 0 2
785 407
785 357
1 1 3 0 0 8320 0 2 1 0 0 3
789 508
776 508
776 453
0 1 3 0 0 0 0 0 3 65 0 2
305 131
305 85
6 1 5 0 0 8320 0 5 10 0 0 3
809 309
854 309
854 200
2 1 6 0 0 4224 0 4 5 0 0 3
693 272
785 272
785 282
1 0 2 0 0 0 0 6 0 0 8 2
753 327
753 327
2 3 2 0 0 8192 0 5 5 0 0 4
761 309
753 309
753 327
761 327
12 1 7 0 0 4224 0 25 4 0 0 2
635 272
657 272
10 4 8 0 0 8320 0 9 26 0 0 3
583 134
583 137
626 137
11 3 9 0 0 4224 0 9 26 0 0 3
583 143
632 143
632 137
12 2 10 0 0 4224 0 9 26 0 0 3
583 152
638 152
638 137
13 1 11 0 0 4224 0 9 26 0 0 3
583 161
644 161
644 137
1 4 12 0 0 4224 0 7 9 0 0 2
506 134
519 134
1 0 2 0 0 0 0 9 0 0 16 3
519 107
513 107
513 116
2 0 2 0 0 0 0 9 0 0 17 3
519 116
512 116
512 125
3 0 2 0 0 0 0 9 0 0 18 3
519 125
512 125
512 143
5 0 2 0 0 0 0 9 0 0 19 3
519 143
512 143
512 152
6 1 2 0 0 8320 0 9 8 0 0 3
519 152
512 152
512 188
7 0 13 0 0 4096 0 9 0 0 62 2
519 161
483 161
8 0 14 0 0 4096 0 9 0 0 64 2
519 170
430 170
1 9 2 0 0 0 0 8 9 0 0 2
512 188
519 188
10 4 15 0 0 8320 0 15 12 0 0 3
697 363
717 363
717 179
11 3 16 0 0 8320 0 15 12 0 0 3
697 372
723 372
723 179
12 2 17 0 0 8320 0 15 12 0 0 3
697 381
729 381
729 179
13 1 18 0 0 8320 0 15 12 0 0 3
697 390
735 390
735 179
1 0 2 0 0 0 0 11 0 0 29 2
680 190
680 190
0 2 2 0 0 0 0 0 13 29 0 3
686 190
692 190
692 179
4 3 2 0 0 0 0 13 13 0 0 4
680 179
680 190
686 190
686 179
14 1 19 0 0 8320 0 15 13 0 0 4
697 417
706 417
706 179
698 179
0 0 2 0 0 0 0 0 0 32 33 2
618 399
618 417
8 5 2 0 0 0 0 15 15 0 0 4
633 399
618 399
618 372
633 372
9 1 2 0 0 0 0 15 14 0 0 2
633 417
613 417
7 0 20 0 0 4096 0 15 0 0 35 2
633 390
627 390
14 6 20 0 0 8320 0 20 15 0 0 6
638 533
673 533
673 445
627 445
627 381
633 381
4 0 21 0 0 4096 0 15 0 0 52 2
633 363
571 363
3 0 22 0 0 4096 0 15 0 0 53 2
633 354
564 354
2 0 23 0 0 4096 0 15 0 0 54 2
633 345
558 345
1 0 24 0 0 4096 0 15 0 0 55 2
633 336
552 336
1 0 2 0 0 0 0 16 0 0 50 2
642 488
642 488
1 0 2 0 0 0 0 17 0 0 56 2
641 245
641 245
1 0 2 0 0 0 0 18 0 0 44 2
559 524
559 524
1 0 25 0 0 0 0 19 0 0 45 2
568 506
568 506
7 6 2 0 0 0 0 20 20 0 0 4
574 524
559 524
559 515
574 515
8 5 25 0 0 8320 0 20 20 0 0 4
574 533
568 533
568 506
574 506
0 4 21 0 0 4096 0 0 20 52 0 3
571 419
571 497
574 497
0 3 22 0 0 4096 0 0 20 53 0 3
564 401
564 488
574 488
0 2 23 0 0 4096 0 0 20 54 0 3
558 383
558 479
574 479
0 1 24 0 0 4224 0 0 20 55 0 3
550 365
550 470
574 470
9 11 2 0 0 0 0 20 20 0 0 4
638 470
642 470
642 488
638 488
10 1 26 0 0 4224 0 20 21 0 0 2
638 479
647 479
14 8 21 0 0 8320 0 33 25 0 0 3
547 419
571 419
571 290
13 7 22 0 0 8320 0 33 25 0 0 4
547 401
564 401
564 281
571 281
12 6 23 0 0 8320 0 33 25 0 0 4
547 383
558 383
558 272
571 272
11 5 24 0 0 0 0 33 25 0 0 4
547 365
552 365
552 263
571 263
9 11 2 0 0 0 0 25 25 0 0 4
635 227
641 227
641 245
635 245
10 1 27 0 0 4224 0 25 22 0 0 2
635 236
646 236
2 1 2 0 0 0 0 25 24 0 0 2
571 236
541 236
3 0 28 0 0 4096 0 25 0 0 60 2
571 245
559 245
4 0 28 0 0 8320 0 25 0 0 61 3
571 254
559 254
559 227
1 1 28 0 0 0 0 23 25 0 0 2
557 227
571 227
6 1 13 0 0 8320 0 29 33 0 0 3
415 139
483 139
483 347
1 0 14 0 0 0 0 35 0 0 64 2
367 252
335 252
7 1 14 0 0 16512 0 29 34 0 0 6
415 148
430 148
430 226
335 226
335 455
367 455
3 4 3 0 0 0 0 27 29 0 0 4
279 131
305 131
305 157
345 157
2 0 2 0 0 0 0 29 0 0 67 2
351 139
337 139
0 1 2 0 0 0 0 0 29 68 0 3
337 148
337 130
351 130
1 3 2 0 0 0 0 28 29 0 0 3
337 173
337 148
345 148
1 10 2 0 0 0 0 30 34 0 0 2
361 551
361 536
10 1 2 0 0 0 0 35 31 0 0 2
361 333
361 347
4 2 29 0 0 12416 0 36 34 0 0 5
210 548
210 574
307 574
307 464
367 464
3 4 30 0 0 12416 0 36 34 0 0 5
216 548
216 565
298 565
298 482
367 482
2 6 31 0 0 16512 0 36 34 0 0 5
222 548
222 556
289 556
289 500
367 500
1 8 32 0 0 12416 0 36 34 0 0 4
228 548
281 548
281 518
367 518
4 3 33 0 0 16512 0 37 34 0 0 5
209 444
209 463
274 463
274 473
367 473
3 5 34 0 0 16512 0 37 34 0 0 5
215 444
215 456
266 456
266 491
367 491
2 7 35 0 0 16512 0 37 34 0 0 5
221 444
221 449
258 449
258 509
367 509
1 9 36 0 0 12416 0 37 34 0 0 4
227 444
251 444
251 527
367 527
4 2 37 0 0 12416 0 38 35 0 0 5
210 346
210 367
307 367
307 261
367 261
3 4 38 0 0 8320 0 38 35 0 0 5
216 346
216 359
300 359
300 279
367 279
2 6 39 0 0 16512 0 38 35 0 0 5
222 346
222 352
292 352
292 297
367 297
1 8 40 0 0 12416 0 38 35 0 0 4
228 346
284 346
284 315
367 315
4 3 41 0 0 16512 0 39 35 0 0 5
211 246
211 261
276 261
276 270
367 270
3 5 42 0 0 16512 0 39 35 0 0 5
217 246
217 255
267 255
267 288
367 288
2 7 43 0 0 16512 0 39 35 0 0 5
223 246
223 250
259 250
259 306
367 306
1 9 44 0 0 12416 0 39 35 0 0 4
229 246
252 246
252 324
367 324
10 1 2 0 0 0 0 33 32 0 0 3
477 428
477 444
487 444
14 8 45 0 0 8320 0 34 33 0 0 4
431 527
472 527
472 410
483 410
13 6 46 0 0 8320 0 34 33 0 0 4
431 509
465 509
465 392
483 392
12 4 47 0 0 8320 0 34 33 0 0 4
431 491
459 491
459 374
483 374
11 2 48 0 0 8320 0 34 33 0 0 4
431 473
454 473
454 356
483 356
11 3 49 0 0 8320 0 35 33 0 0 4
431 270
448 270
448 365
483 365
12 5 50 0 0 8320 0 35 33 0 0 4
431 288
443 288
443 383
483 383
13 7 51 0 0 8320 0 35 33 0 0 4
431 306
437 306
437 401
483 401
14 9 52 0 0 4224 0 35 33 0 0 3
431 324
431 419
483 419
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
