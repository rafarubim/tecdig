CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 100 10
176 80 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 692 69 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43232.7 0
0
9 Inverter~
13 272 642 0 2 22
0 4 5
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4F
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
391 0 0
2
43232.7 0
0
9 2-In AND~
219 181 603 0 3 22
0 3 5 6
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U8A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3124 0 0
2
43232.7 0
0
8 2-In OR~
219 345 203 0 3 22
0 4 9 8
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U7C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3421 0 0
2
43232.7 0
0
9 Inverter~
13 284 180 0 2 22
0 7 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
8157 0 0
2
43232.7 0
0
8 2-In OR~
219 431 536 0 3 22
0 4 10 11
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U7B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5572 0 0
2
43232.7 0
0
9 Inverter~
13 186 407 0 2 22
0 3 13
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U4D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
8901 0 0
2
43232.7 0
0
8 2-In OR~
219 186 530 0 3 22
0 6 14 3
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U7A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7361 0 0
2
43232.7 0
0
9 2-In AND~
219 262 321 0 3 22
0 12 13 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4747 0 0
2
43232.7 0
0
9 2-In AND~
219 631 422 0 3 22
0 17 16 14
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
972 0 0
2
43232.7 0
0
9 Inverter~
13 312 321 0 2 22
0 15 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3472 0 0
2
43232.7 0
0
7 Ground~
168 362 414 0 1 3
0 2
0
0 0 53360 270
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9998 0 0
2
43232.7 0
0
9 2-In AND~
219 559 421 0 3 22
0 19 20 10
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3536 0 0
2
43232.7 0
0
9 Inverter~
13 422 377 0 2 22
0 20 22
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
4597 0 0
2
43232.7 0
0
9 2-In AND~
219 385 386 0 3 22
0 19 22 21
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U6A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3835 0 0
2
43232.7 0
0
14 Logic Display~
6 475 484 0 1 2
10 23
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
43232.7 0
0
5 4013~
219 383 485 0 6 22
0 2 21 12 11 26 23
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
5616 0 0
2
43232.7 0
0
7 Ground~
168 509 249 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9323 0 0
2
43232.7 0
0
7 74LS290
153 387 303 0 10 21
0 2 2 8 8 18 16 20 24 25
16
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 0 0 0 0
1 U
317 0 0
2
43232.7 7
0
7 74LS290
153 551 304 0 10 21
0 2 2 8 8 20 19 27 28 17
19
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 512 0 0 0 0
1 U
3108 0 0
2
43232.7 6
0
12 Hex Display~
7 469 164 0 18 19
10 16 25 24 20 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4299 0 0
2
43232.7 5
0
12 Hex Display~
7 420 164 0 16 19
10 19 17 29 30 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
9672 0 0
2
43232.7 4
0
7 Pulser~
4 105 321 0 10 12
0 31 32 12 33 0 0 10 10 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7876 0 0
2
43232.7 3
0
5 4071~
219 210 213 0 3 22
0 7 12 7
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
6369 0 0
2
43232.7 2
0
7 Ground~
168 292 284 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9172 0 0
2
43232.7 0
0
46
1 0 3 0 0 12416 0 3 0 0 5 5
171 624
171 642
148 642
148 467
189 467
1 0 4 0 0 4096 0 2 0 0 7 3
293 642
475 642
475 545
2 2 5 0 0 8320 0 3 2 0 0 3
189 624
189 642
257 642
3 1 6 0 0 4224 0 3 8 0 0 2
180 579
180 546
1 3 3 0 0 0 0 7 8 0 0 2
189 425
189 500
3 0 7 0 0 8192 0 24 0 0 14 3
243 213
259 213
259 180
1 0 4 0 0 8320 0 6 0 0 8 3
450 545
692 545
692 108
1 1 4 0 0 0 0 4 1 0 0 4
357 187
357 108
692 108
692 81
3 0 8 0 0 4096 0 20 0 0 10 2
519 295
494 295
4 0 8 0 0 12416 0 20 0 0 12 4
519 304
494 304
494 243
348 243
3 0 8 0 0 0 0 19 0 0 12 2
355 294
348 294
3 4 8 0 0 0 0 4 19 0 0 3
348 233
348 303
355 303
2 2 9 0 0 4224 0 5 4 0 0 3
305 180
339 180
339 187
1 1 7 0 0 4224 0 5 24 0 0 4
269 180
189 180
189 204
197 204
2 3 10 0 0 4224 0 6 13 0 0 3
450 527
557 527
557 444
4 3 11 0 0 4224 0 17 6 0 0 3
383 491
383 536
404 536
3 0 12 0 0 8320 0 17 0 0 21 3
359 467
213 467
213 312
2 2 13 0 0 8320 0 9 7 0 0 3
238 330
189 330
189 389
2 3 14 0 0 8320 0 8 10 0 0 4
198 546
198 573
629 573
629 445
2 0 12 0 0 0 0 24 0 0 21 3
197 222
189 222
189 312
3 1 12 0 0 0 0 23 9 0 0 2
129 312
238 312
3 1 15 0 0 12416 0 9 11 0 0 4
283 321
282 321
282 321
297 321
2 0 16 0 0 8320 0 10 0 0 42 5
620 400
620 362
478 362
478 345
434 345
1 0 17 0 0 4096 0 10 0 0 35 3
638 400
638 351
590 351
2 5 18 0 0 4224 0 11 19 0 0 2
333 321
349 321
1 1 2 0 0 8320 0 17 12 0 0 3
383 428
383 415
369 415
1 0 19 0 0 8192 0 13 0 0 32 3
566 399
566 395
508 395
2 0 20 0 0 8192 0 13 0 0 29 3
548 399
548 377
459 377
1 0 20 0 0 8320 0 14 0 0 38 3
443 377
460 377
460 276
2 3 21 0 0 8320 0 17 15 0 0 4
359 449
340 449
340 386
358 386
2 2 22 0 0 4224 0 15 14 0 0 2
403 377
407 377
1 0 19 0 0 4096 0 15 0 0 34 3
403 395
509 395
509 345
6 1 23 0 0 4224 0 17 16 0 0 3
407 449
475 449
475 470
6 0 19 0 0 0 0 20 0 0 39 5
513 331
509 331
509 345
587 345
587 331
2 9 17 0 0 8320 0 22 20 0 0 5
423 188
423 351
591 351
591 313
583 313
1 0 2 0 0 0 0 20 0 0 37 2
519 277
509 277
1 2 2 0 0 4096 0 18 20 0 0 3
509 257
509 286
519 286
5 0 20 0 0 0 0 20 0 0 43 4
513 322
486 322
486 276
460 276
10 1 19 0 0 12416 0 20 22 0 0 5
583 331
587 331
587 196
429 196
429 188
1 0 2 0 0 4096 0 19 0 0 41 3
355 276
316 276
316 285
2 1 2 0 0 4224 0 19 25 0 0 2
355 285
299 285
6 0 16 0 0 0 0 19 0 0 46 5
349 330
340 330
340 345
435 345
435 330
7 4 20 0 0 128 0 19 21 0 0 3
419 276
460 276
460 188
8 3 24 0 0 8320 0 19 21 0 0 3
419 294
466 294
466 188
9 2 25 0 0 8320 0 19 21 0 0 3
419 312
472 312
472 188
10 1 16 0 0 128 0 19 21 0 0 3
419 330
478 330
478 188
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
