CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 21 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 F:\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
176 550 1918 1019
9437202 0
0
6 Title:
5 Name:
0
0
0
8
12 Hex Display~
7 649 545 0 16 19
10 11 10 9 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4747 0 0
2
5.89841e-315 0
0
12 Hex Display~
7 608 546 0 16 19
10 7 6 5 4 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.89841e-315 0
0
9 2-In AND~
219 636 461 0 3 22
0 10 11 12
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
5.89841e-315 0
0
7 Ground~
168 697 322 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
5.89841e-315 0
0
7 74LS290
153 729 385 0 10 21
0 2 2 6 12 8 7 4 5 6
7
0
0 0 4336 0
7 74LS290
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.89841e-315 0
0
7 Ground~
168 561 320 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89841e-315 0
0
7 74LS290
153 593 384 0 10 21
0 2 2 6 12 3 11 8 9 10
11
0
0 0 4336 0
7 74LS290
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.89841e-315 0
0
7 Pulser~
4 467 411 0 10 12
0 13 14 3 15 0 0 30 30 31
7
0
0 0 4144 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
5.89841e-315 0
0
22
3 5 3 0 0 4224 0 8 7 0 0 2
491 402
555 402
7 4 4 0 0 8320 0 5 2 0 0 5
761 358
790 358
790 608
599 608
599 570
8 3 5 0 0 8320 0 5 2 0 0 5
761 376
783 376
783 603
605 603
605 570
0 2 6 0 0 8192 0 0 2 13 0 4
776 492
776 597
611 597
611 570
0 1 7 0 0 4224 0 0 2 19 0 4
761 430
761 592
617 592
617 570
0 4 8 0 0 12416 0 0 1 18 0 6
667 403
667 465
706 465
706 586
640 586
640 569
8 3 9 0 0 24704 0 7 1 0 0 9
625 375
648 375
648 421
662 421
662 470
701 470
701 579
646 579
646 569
0 2 10 0 0 16512 0 0 1 14 0 7
643 425
658 425
658 474
697 474
697 573
652 573
652 569
0 1 11 0 0 16512 0 0 1 15 0 6
625 430
655 430
655 478
693 478
693 569
658 569
3 4 12 0 0 8320 0 3 7 0 0 4
634 484
550 484
550 384
561 384
3 4 12 0 0 0 0 3 5 0 0 4
634 484
685 484
685 385
697 385
3 0 6 0 0 0 0 5 0 0 13 3
697 376
677 376
677 493
9 3 6 0 0 12416 0 5 7 0 0 6
761 394
776 394
776 493
542 493
542 375
561 375
1 9 10 0 0 0 0 3 7 0 0 3
643 439
643 393
625 393
2 0 11 0 0 0 0 3 0 0 20 2
625 439
625 430
1 1 2 0 0 4096 0 5 4 0 0 2
697 358
697 330
2 1 2 0 0 0 0 5 5 0 0 2
697 367
697 358
7 5 8 0 0 0 0 7 5 0 0 4
625 357
658 357
658 403
691 403
6 10 7 0 0 0 0 5 5 0 0 4
691 412
691 430
761 430
761 412
6 10 11 0 0 0 0 7 7 0 0 4
555 411
555 430
625 430
625 411
1 1 2 0 0 4224 0 7 6 0 0 2
561 357
561 328
2 1 2 0 0 0 0 7 7 0 0 2
561 366
561 357
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
